
    wire dl_reset;
    wire dl_clock;
    assign dl_reset = ap_rst_n;
    assign dl_clock = ap_clk;
    wire [2:0] proc_0_data_FIFO_blk;
    wire [2:0] proc_0_data_PIPO_blk;
    wire [2:0] proc_0_start_FIFO_blk;
    wire [2:0] proc_0_TLF_FIFO_blk;
    wire [2:0] proc_0_input_sync_blk;
    wire [2:0] proc_0_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_0;
    reg [2:0] proc_dep_vld_vec_0_reg;
    wire [2:0] in_chan_dep_vld_vec_0;
    wire [77:0] in_chan_dep_data_vec_0;
    wire [2:0] token_in_vec_0;
    wire [2:0] out_chan_dep_vld_vec_0;
    wire [25:0] out_chan_dep_data_0;
    wire [2:0] token_out_vec_0;
    wire dl_detect_out_0;
    wire dep_chan_vld_1_0;
    wire [25:0] dep_chan_data_1_0;
    wire token_1_0;
    wire dep_chan_vld_2_0;
    wire [25:0] dep_chan_data_2_0;
    wire token_2_0;
    wire dep_chan_vld_25_0;
    wire [25:0] dep_chan_data_25_0;
    wire token_25_0;
    wire [3:0] proc_1_data_FIFO_blk;
    wire [3:0] proc_1_data_PIPO_blk;
    wire [3:0] proc_1_start_FIFO_blk;
    wire [3:0] proc_1_TLF_FIFO_blk;
    wire [3:0] proc_1_input_sync_blk;
    wire [3:0] proc_1_output_sync_blk;
    wire [3:0] proc_dep_vld_vec_1;
    reg [3:0] proc_dep_vld_vec_1_reg;
    wire [3:0] in_chan_dep_vld_vec_1;
    wire [103:0] in_chan_dep_data_vec_1;
    wire [3:0] token_in_vec_1;
    wire [3:0] out_chan_dep_vld_vec_1;
    wire [25:0] out_chan_dep_data_1;
    wire [3:0] token_out_vec_1;
    wire dl_detect_out_1;
    wire dep_chan_vld_0_1;
    wire [25:0] dep_chan_data_0_1;
    wire token_0_1;
    wire dep_chan_vld_2_1;
    wire [25:0] dep_chan_data_2_1;
    wire token_2_1;
    wire dep_chan_vld_3_1;
    wire [25:0] dep_chan_data_3_1;
    wire token_3_1;
    wire dep_chan_vld_4_1;
    wire [25:0] dep_chan_data_4_1;
    wire token_4_1;
    wire [3:0] proc_2_data_FIFO_blk;
    wire [3:0] proc_2_data_PIPO_blk;
    wire [3:0] proc_2_start_FIFO_blk;
    wire [3:0] proc_2_TLF_FIFO_blk;
    wire [3:0] proc_2_input_sync_blk;
    wire [3:0] proc_2_output_sync_blk;
    wire [3:0] proc_dep_vld_vec_2;
    reg [3:0] proc_dep_vld_vec_2_reg;
    wire [3:0] in_chan_dep_vld_vec_2;
    wire [103:0] in_chan_dep_data_vec_2;
    wire [3:0] token_in_vec_2;
    wire [3:0] out_chan_dep_vld_vec_2;
    wire [25:0] out_chan_dep_data_2;
    wire [3:0] token_out_vec_2;
    wire dl_detect_out_2;
    wire dep_chan_vld_0_2;
    wire [25:0] dep_chan_data_0_2;
    wire token_0_2;
    wire dep_chan_vld_1_2;
    wire [25:0] dep_chan_data_1_2;
    wire token_1_2;
    wire dep_chan_vld_3_2;
    wire [25:0] dep_chan_data_3_2;
    wire token_3_2;
    wire dep_chan_vld_20_2;
    wire [25:0] dep_chan_data_20_2;
    wire token_20_2;
    wire [2:0] proc_3_data_FIFO_blk;
    wire [2:0] proc_3_data_PIPO_blk;
    wire [2:0] proc_3_start_FIFO_blk;
    wire [2:0] proc_3_TLF_FIFO_blk;
    wire [2:0] proc_3_input_sync_blk;
    wire [2:0] proc_3_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_3;
    reg [2:0] proc_dep_vld_vec_3_reg;
    wire [2:0] in_chan_dep_vld_vec_3;
    wire [77:0] in_chan_dep_data_vec_3;
    wire [2:0] token_in_vec_3;
    wire [2:0] out_chan_dep_vld_vec_3;
    wire [25:0] out_chan_dep_data_3;
    wire [2:0] token_out_vec_3;
    wire dl_detect_out_3;
    wire dep_chan_vld_1_3;
    wire [25:0] dep_chan_data_1_3;
    wire token_1_3;
    wire dep_chan_vld_2_3;
    wire [25:0] dep_chan_data_2_3;
    wire token_2_3;
    wire dep_chan_vld_25_3;
    wire [25:0] dep_chan_data_25_3;
    wire token_25_3;
    wire [1:0] proc_4_data_FIFO_blk;
    wire [1:0] proc_4_data_PIPO_blk;
    wire [1:0] proc_4_start_FIFO_blk;
    wire [1:0] proc_4_TLF_FIFO_blk;
    wire [1:0] proc_4_input_sync_blk;
    wire [1:0] proc_4_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_4;
    reg [1:0] proc_dep_vld_vec_4_reg;
    wire [1:0] in_chan_dep_vld_vec_4;
    wire [51:0] in_chan_dep_data_vec_4;
    wire [1:0] token_in_vec_4;
    wire [1:0] out_chan_dep_vld_vec_4;
    wire [25:0] out_chan_dep_data_4;
    wire [1:0] token_out_vec_4;
    wire dl_detect_out_4;
    wire dep_chan_vld_1_4;
    wire [25:0] dep_chan_data_1_4;
    wire token_1_4;
    wire dep_chan_vld_5_4;
    wire [25:0] dep_chan_data_5_4;
    wire token_5_4;
    wire [1:0] proc_5_data_FIFO_blk;
    wire [1:0] proc_5_data_PIPO_blk;
    wire [1:0] proc_5_start_FIFO_blk;
    wire [1:0] proc_5_TLF_FIFO_blk;
    wire [1:0] proc_5_input_sync_blk;
    wire [1:0] proc_5_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_5;
    reg [1:0] proc_dep_vld_vec_5_reg;
    wire [1:0] in_chan_dep_vld_vec_5;
    wire [51:0] in_chan_dep_data_vec_5;
    wire [1:0] token_in_vec_5;
    wire [1:0] out_chan_dep_vld_vec_5;
    wire [25:0] out_chan_dep_data_5;
    wire [1:0] token_out_vec_5;
    wire dl_detect_out_5;
    wire dep_chan_vld_4_5;
    wire [25:0] dep_chan_data_4_5;
    wire token_4_5;
    wire dep_chan_vld_6_5;
    wire [25:0] dep_chan_data_6_5;
    wire token_6_5;
    wire [2:0] proc_6_data_FIFO_blk;
    wire [2:0] proc_6_data_PIPO_blk;
    wire [2:0] proc_6_start_FIFO_blk;
    wire [2:0] proc_6_TLF_FIFO_blk;
    wire [2:0] proc_6_input_sync_blk;
    wire [2:0] proc_6_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_6;
    reg [2:0] proc_dep_vld_vec_6_reg;
    wire [2:0] in_chan_dep_vld_vec_6;
    wire [77:0] in_chan_dep_data_vec_6;
    wire [2:0] token_in_vec_6;
    wire [2:0] out_chan_dep_vld_vec_6;
    wire [25:0] out_chan_dep_data_6;
    wire [2:0] token_out_vec_6;
    wire dl_detect_out_6;
    wire dep_chan_vld_5_6;
    wire [25:0] dep_chan_data_5_6;
    wire token_5_6;
    wire dep_chan_vld_7_6;
    wire [25:0] dep_chan_data_7_6;
    wire token_7_6;
    wire dep_chan_vld_8_6;
    wire [25:0] dep_chan_data_8_6;
    wire token_8_6;
    wire [1:0] proc_7_data_FIFO_blk;
    wire [1:0] proc_7_data_PIPO_blk;
    wire [1:0] proc_7_start_FIFO_blk;
    wire [1:0] proc_7_TLF_FIFO_blk;
    wire [1:0] proc_7_input_sync_blk;
    wire [1:0] proc_7_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_7;
    reg [1:0] proc_dep_vld_vec_7_reg;
    wire [1:0] in_chan_dep_vld_vec_7;
    wire [51:0] in_chan_dep_data_vec_7;
    wire [1:0] token_in_vec_7;
    wire [1:0] out_chan_dep_vld_vec_7;
    wire [25:0] out_chan_dep_data_7;
    wire [1:0] token_out_vec_7;
    wire dl_detect_out_7;
    wire dep_chan_vld_6_7;
    wire [25:0] dep_chan_data_6_7;
    wire token_6_7;
    wire dep_chan_vld_9_7;
    wire [25:0] dep_chan_data_9_7;
    wire token_9_7;
    wire [1:0] proc_8_data_FIFO_blk;
    wire [1:0] proc_8_data_PIPO_blk;
    wire [1:0] proc_8_start_FIFO_blk;
    wire [1:0] proc_8_TLF_FIFO_blk;
    wire [1:0] proc_8_input_sync_blk;
    wire [1:0] proc_8_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_8;
    reg [1:0] proc_dep_vld_vec_8_reg;
    wire [1:0] in_chan_dep_vld_vec_8;
    wire [51:0] in_chan_dep_data_vec_8;
    wire [1:0] token_in_vec_8;
    wire [1:0] out_chan_dep_vld_vec_8;
    wire [25:0] out_chan_dep_data_8;
    wire [1:0] token_out_vec_8;
    wire dl_detect_out_8;
    wire dep_chan_vld_6_8;
    wire [25:0] dep_chan_data_6_8;
    wire token_6_8;
    wire dep_chan_vld_11_8;
    wire [25:0] dep_chan_data_11_8;
    wire token_11_8;
    wire [1:0] proc_9_data_FIFO_blk;
    wire [1:0] proc_9_data_PIPO_blk;
    wire [1:0] proc_9_start_FIFO_blk;
    wire [1:0] proc_9_TLF_FIFO_blk;
    wire [1:0] proc_9_input_sync_blk;
    wire [1:0] proc_9_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_9;
    reg [1:0] proc_dep_vld_vec_9_reg;
    wire [1:0] in_chan_dep_vld_vec_9;
    wire [51:0] in_chan_dep_data_vec_9;
    wire [1:0] token_in_vec_9;
    wire [1:0] out_chan_dep_vld_vec_9;
    wire [25:0] out_chan_dep_data_9;
    wire [1:0] token_out_vec_9;
    wire dl_detect_out_9;
    wire dep_chan_vld_7_9;
    wire [25:0] dep_chan_data_7_9;
    wire token_7_9;
    wire dep_chan_vld_10_9;
    wire [25:0] dep_chan_data_10_9;
    wire token_10_9;
    wire [2:0] proc_10_data_FIFO_blk;
    wire [2:0] proc_10_data_PIPO_blk;
    wire [2:0] proc_10_start_FIFO_blk;
    wire [2:0] proc_10_TLF_FIFO_blk;
    wire [2:0] proc_10_input_sync_blk;
    wire [2:0] proc_10_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_10;
    reg [2:0] proc_dep_vld_vec_10_reg;
    wire [2:0] in_chan_dep_vld_vec_10;
    wire [77:0] in_chan_dep_data_vec_10;
    wire [2:0] token_in_vec_10;
    wire [2:0] out_chan_dep_vld_vec_10;
    wire [25:0] out_chan_dep_data_10;
    wire [2:0] token_out_vec_10;
    wire dl_detect_out_10;
    wire dep_chan_vld_9_10;
    wire [25:0] dep_chan_data_9_10;
    wire token_9_10;
    wire dep_chan_vld_13_10;
    wire [25:0] dep_chan_data_13_10;
    wire token_13_10;
    wire dep_chan_vld_18_10;
    wire [25:0] dep_chan_data_18_10;
    wire token_18_10;
    wire [1:0] proc_11_data_FIFO_blk;
    wire [1:0] proc_11_data_PIPO_blk;
    wire [1:0] proc_11_start_FIFO_blk;
    wire [1:0] proc_11_TLF_FIFO_blk;
    wire [1:0] proc_11_input_sync_blk;
    wire [1:0] proc_11_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_11;
    reg [1:0] proc_dep_vld_vec_11_reg;
    wire [1:0] in_chan_dep_vld_vec_11;
    wire [51:0] in_chan_dep_data_vec_11;
    wire [1:0] token_in_vec_11;
    wire [1:0] out_chan_dep_vld_vec_11;
    wire [25:0] out_chan_dep_data_11;
    wire [1:0] token_out_vec_11;
    wire dl_detect_out_11;
    wire dep_chan_vld_8_11;
    wire [25:0] dep_chan_data_8_11;
    wire token_8_11;
    wire dep_chan_vld_12_11;
    wire [25:0] dep_chan_data_12_11;
    wire token_12_11;
    wire [1:0] proc_12_data_FIFO_blk;
    wire [1:0] proc_12_data_PIPO_blk;
    wire [1:0] proc_12_start_FIFO_blk;
    wire [1:0] proc_12_TLF_FIFO_blk;
    wire [1:0] proc_12_input_sync_blk;
    wire [1:0] proc_12_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_12;
    reg [1:0] proc_dep_vld_vec_12_reg;
    wire [1:0] in_chan_dep_vld_vec_12;
    wire [51:0] in_chan_dep_data_vec_12;
    wire [1:0] token_in_vec_12;
    wire [1:0] out_chan_dep_vld_vec_12;
    wire [25:0] out_chan_dep_data_12;
    wire [1:0] token_out_vec_12;
    wire dl_detect_out_12;
    wire dep_chan_vld_11_12;
    wire [25:0] dep_chan_data_11_12;
    wire token_11_12;
    wire dep_chan_vld_14_12;
    wire [25:0] dep_chan_data_14_12;
    wire token_14_12;
    wire [1:0] proc_13_data_FIFO_blk;
    wire [1:0] proc_13_data_PIPO_blk;
    wire [1:0] proc_13_start_FIFO_blk;
    wire [1:0] proc_13_TLF_FIFO_blk;
    wire [1:0] proc_13_input_sync_blk;
    wire [1:0] proc_13_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_13;
    reg [1:0] proc_dep_vld_vec_13_reg;
    wire [1:0] in_chan_dep_vld_vec_13;
    wire [51:0] in_chan_dep_data_vec_13;
    wire [1:0] token_in_vec_13;
    wire [1:0] out_chan_dep_vld_vec_13;
    wire [25:0] out_chan_dep_data_13;
    wire [1:0] token_out_vec_13;
    wire dl_detect_out_13;
    wire dep_chan_vld_10_13;
    wire [25:0] dep_chan_data_10_13;
    wire token_10_13;
    wire dep_chan_vld_15_13;
    wire [25:0] dep_chan_data_15_13;
    wire token_15_13;
    wire [1:0] proc_14_data_FIFO_blk;
    wire [1:0] proc_14_data_PIPO_blk;
    wire [1:0] proc_14_start_FIFO_blk;
    wire [1:0] proc_14_TLF_FIFO_blk;
    wire [1:0] proc_14_input_sync_blk;
    wire [1:0] proc_14_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_14;
    reg [1:0] proc_dep_vld_vec_14_reg;
    wire [1:0] in_chan_dep_vld_vec_14;
    wire [51:0] in_chan_dep_data_vec_14;
    wire [1:0] token_in_vec_14;
    wire [1:0] out_chan_dep_vld_vec_14;
    wire [25:0] out_chan_dep_data_14;
    wire [1:0] token_out_vec_14;
    wire dl_detect_out_14;
    wire dep_chan_vld_12_14;
    wire [25:0] dep_chan_data_12_14;
    wire token_12_14;
    wire dep_chan_vld_16_14;
    wire [25:0] dep_chan_data_16_14;
    wire token_16_14;
    wire [1:0] proc_15_data_FIFO_blk;
    wire [1:0] proc_15_data_PIPO_blk;
    wire [1:0] proc_15_start_FIFO_blk;
    wire [1:0] proc_15_TLF_FIFO_blk;
    wire [1:0] proc_15_input_sync_blk;
    wire [1:0] proc_15_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_15;
    reg [1:0] proc_dep_vld_vec_15_reg;
    wire [1:0] in_chan_dep_vld_vec_15;
    wire [51:0] in_chan_dep_data_vec_15;
    wire [1:0] token_in_vec_15;
    wire [1:0] out_chan_dep_vld_vec_15;
    wire [25:0] out_chan_dep_data_15;
    wire [1:0] token_out_vec_15;
    wire dl_detect_out_15;
    wire dep_chan_vld_13_15;
    wire [25:0] dep_chan_data_13_15;
    wire token_13_15;
    wire dep_chan_vld_16_15;
    wire [25:0] dep_chan_data_16_15;
    wire token_16_15;
    wire [2:0] proc_16_data_FIFO_blk;
    wire [2:0] proc_16_data_PIPO_blk;
    wire [2:0] proc_16_start_FIFO_blk;
    wire [2:0] proc_16_TLF_FIFO_blk;
    wire [2:0] proc_16_input_sync_blk;
    wire [2:0] proc_16_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_16;
    reg [2:0] proc_dep_vld_vec_16_reg;
    wire [2:0] in_chan_dep_vld_vec_16;
    wire [77:0] in_chan_dep_data_vec_16;
    wire [2:0] token_in_vec_16;
    wire [2:0] out_chan_dep_vld_vec_16;
    wire [25:0] out_chan_dep_data_16;
    wire [2:0] token_out_vec_16;
    wire dl_detect_out_16;
    wire dep_chan_vld_14_16;
    wire [25:0] dep_chan_data_14_16;
    wire token_14_16;
    wire dep_chan_vld_15_16;
    wire [25:0] dep_chan_data_15_16;
    wire token_15_16;
    wire dep_chan_vld_17_16;
    wire [25:0] dep_chan_data_17_16;
    wire token_17_16;
    wire [1:0] proc_17_data_FIFO_blk;
    wire [1:0] proc_17_data_PIPO_blk;
    wire [1:0] proc_17_start_FIFO_blk;
    wire [1:0] proc_17_TLF_FIFO_blk;
    wire [1:0] proc_17_input_sync_blk;
    wire [1:0] proc_17_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_17;
    reg [1:0] proc_dep_vld_vec_17_reg;
    wire [1:0] in_chan_dep_vld_vec_17;
    wire [51:0] in_chan_dep_data_vec_17;
    wire [1:0] token_in_vec_17;
    wire [1:0] out_chan_dep_vld_vec_17;
    wire [25:0] out_chan_dep_data_17;
    wire [1:0] token_out_vec_17;
    wire dl_detect_out_17;
    wire dep_chan_vld_16_17;
    wire [25:0] dep_chan_data_16_17;
    wire token_16_17;
    wire dep_chan_vld_18_17;
    wire [25:0] dep_chan_data_18_17;
    wire token_18_17;
    wire [2:0] proc_18_data_FIFO_blk;
    wire [2:0] proc_18_data_PIPO_blk;
    wire [2:0] proc_18_start_FIFO_blk;
    wire [2:0] proc_18_TLF_FIFO_blk;
    wire [2:0] proc_18_input_sync_blk;
    wire [2:0] proc_18_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_18;
    reg [2:0] proc_dep_vld_vec_18_reg;
    wire [2:0] in_chan_dep_vld_vec_18;
    wire [77:0] in_chan_dep_data_vec_18;
    wire [2:0] token_in_vec_18;
    wire [2:0] out_chan_dep_vld_vec_18;
    wire [25:0] out_chan_dep_data_18;
    wire [2:0] token_out_vec_18;
    wire dl_detect_out_18;
    wire dep_chan_vld_10_18;
    wire [25:0] dep_chan_data_10_18;
    wire token_10_18;
    wire dep_chan_vld_17_18;
    wire [25:0] dep_chan_data_17_18;
    wire token_17_18;
    wire dep_chan_vld_19_18;
    wire [25:0] dep_chan_data_19_18;
    wire token_19_18;
    wire [1:0] proc_19_data_FIFO_blk;
    wire [1:0] proc_19_data_PIPO_blk;
    wire [1:0] proc_19_start_FIFO_blk;
    wire [1:0] proc_19_TLF_FIFO_blk;
    wire [1:0] proc_19_input_sync_blk;
    wire [1:0] proc_19_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_19;
    reg [1:0] proc_dep_vld_vec_19_reg;
    wire [1:0] in_chan_dep_vld_vec_19;
    wire [51:0] in_chan_dep_data_vec_19;
    wire [1:0] token_in_vec_19;
    wire [1:0] out_chan_dep_vld_vec_19;
    wire [25:0] out_chan_dep_data_19;
    wire [1:0] token_out_vec_19;
    wire dl_detect_out_19;
    wire dep_chan_vld_18_19;
    wire [25:0] dep_chan_data_18_19;
    wire token_18_19;
    wire dep_chan_vld_20_19;
    wire [25:0] dep_chan_data_20_19;
    wire token_20_19;
    wire [2:0] proc_20_data_FIFO_blk;
    wire [2:0] proc_20_data_PIPO_blk;
    wire [2:0] proc_20_start_FIFO_blk;
    wire [2:0] proc_20_TLF_FIFO_blk;
    wire [2:0] proc_20_input_sync_blk;
    wire [2:0] proc_20_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_20;
    reg [2:0] proc_dep_vld_vec_20_reg;
    wire [2:0] in_chan_dep_vld_vec_20;
    wire [77:0] in_chan_dep_data_vec_20;
    wire [2:0] token_in_vec_20;
    wire [2:0] out_chan_dep_vld_vec_20;
    wire [25:0] out_chan_dep_data_20;
    wire [2:0] token_out_vec_20;
    wire dl_detect_out_20;
    wire dep_chan_vld_2_20;
    wire [25:0] dep_chan_data_2_20;
    wire token_2_20;
    wire dep_chan_vld_19_20;
    wire [25:0] dep_chan_data_19_20;
    wire token_19_20;
    wire dep_chan_vld_21_20;
    wire [25:0] dep_chan_data_21_20;
    wire token_21_20;
    wire [1:0] proc_21_data_FIFO_blk;
    wire [1:0] proc_21_data_PIPO_blk;
    wire [1:0] proc_21_start_FIFO_blk;
    wire [1:0] proc_21_TLF_FIFO_blk;
    wire [1:0] proc_21_input_sync_blk;
    wire [1:0] proc_21_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_21;
    reg [1:0] proc_dep_vld_vec_21_reg;
    wire [1:0] in_chan_dep_vld_vec_21;
    wire [51:0] in_chan_dep_data_vec_21;
    wire [1:0] token_in_vec_21;
    wire [1:0] out_chan_dep_vld_vec_21;
    wire [25:0] out_chan_dep_data_21;
    wire [1:0] token_out_vec_21;
    wire dl_detect_out_21;
    wire dep_chan_vld_20_21;
    wire [25:0] dep_chan_data_20_21;
    wire token_20_21;
    wire dep_chan_vld_22_21;
    wire [25:0] dep_chan_data_22_21;
    wire token_22_21;
    wire [1:0] proc_22_data_FIFO_blk;
    wire [1:0] proc_22_data_PIPO_blk;
    wire [1:0] proc_22_start_FIFO_blk;
    wire [1:0] proc_22_TLF_FIFO_blk;
    wire [1:0] proc_22_input_sync_blk;
    wire [1:0] proc_22_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_22;
    reg [1:0] proc_dep_vld_vec_22_reg;
    wire [1:0] in_chan_dep_vld_vec_22;
    wire [51:0] in_chan_dep_data_vec_22;
    wire [1:0] token_in_vec_22;
    wire [1:0] out_chan_dep_vld_vec_22;
    wire [25:0] out_chan_dep_data_22;
    wire [1:0] token_out_vec_22;
    wire dl_detect_out_22;
    wire dep_chan_vld_21_22;
    wire [25:0] dep_chan_data_21_22;
    wire token_21_22;
    wire dep_chan_vld_23_22;
    wire [25:0] dep_chan_data_23_22;
    wire token_23_22;
    wire [1:0] proc_23_data_FIFO_blk;
    wire [1:0] proc_23_data_PIPO_blk;
    wire [1:0] proc_23_start_FIFO_blk;
    wire [1:0] proc_23_TLF_FIFO_blk;
    wire [1:0] proc_23_input_sync_blk;
    wire [1:0] proc_23_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_23;
    reg [1:0] proc_dep_vld_vec_23_reg;
    wire [1:0] in_chan_dep_vld_vec_23;
    wire [51:0] in_chan_dep_data_vec_23;
    wire [1:0] token_in_vec_23;
    wire [1:0] out_chan_dep_vld_vec_23;
    wire [25:0] out_chan_dep_data_23;
    wire [1:0] token_out_vec_23;
    wire dl_detect_out_23;
    wire dep_chan_vld_22_23;
    wire [25:0] dep_chan_data_22_23;
    wire token_22_23;
    wire dep_chan_vld_24_23;
    wire [25:0] dep_chan_data_24_23;
    wire token_24_23;
    wire [1:0] proc_24_data_FIFO_blk;
    wire [1:0] proc_24_data_PIPO_blk;
    wire [1:0] proc_24_start_FIFO_blk;
    wire [1:0] proc_24_TLF_FIFO_blk;
    wire [1:0] proc_24_input_sync_blk;
    wire [1:0] proc_24_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_24;
    reg [1:0] proc_dep_vld_vec_24_reg;
    wire [1:0] in_chan_dep_vld_vec_24;
    wire [51:0] in_chan_dep_data_vec_24;
    wire [1:0] token_in_vec_24;
    wire [1:0] out_chan_dep_vld_vec_24;
    wire [25:0] out_chan_dep_data_24;
    wire [1:0] token_out_vec_24;
    wire dl_detect_out_24;
    wire dep_chan_vld_23_24;
    wire [25:0] dep_chan_data_23_24;
    wire token_23_24;
    wire dep_chan_vld_25_24;
    wire [25:0] dep_chan_data_25_24;
    wire token_25_24;
    wire [2:0] proc_25_data_FIFO_blk;
    wire [2:0] proc_25_data_PIPO_blk;
    wire [2:0] proc_25_start_FIFO_blk;
    wire [2:0] proc_25_TLF_FIFO_blk;
    wire [2:0] proc_25_input_sync_blk;
    wire [2:0] proc_25_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_25;
    reg [2:0] proc_dep_vld_vec_25_reg;
    wire [2:0] in_chan_dep_vld_vec_25;
    wire [77:0] in_chan_dep_data_vec_25;
    wire [2:0] token_in_vec_25;
    wire [2:0] out_chan_dep_vld_vec_25;
    wire [25:0] out_chan_dep_data_25;
    wire [2:0] token_out_vec_25;
    wire dl_detect_out_25;
    wire dep_chan_vld_0_25;
    wire [25:0] dep_chan_data_0_25;
    wire token_0_25;
    wire dep_chan_vld_3_25;
    wire [25:0] dep_chan_data_3_25;
    wire token_3_25;
    wire dep_chan_vld_24_25;
    wire [25:0] dep_chan_data_24_25;
    wire token_24_25;
    wire [25:0] dl_in_vec;
    wire dl_detect_out;
    wire token_clear;
    reg [25:0] origin;

reg [15:0] trans_in_cnt_0;// for process Loop_VITIS_LOOP_67_1_proc39_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_0 <= 16'h0;
    end
    else if (Loop_VITIS_LOOP_67_1_proc39_U0.start_write == 1'b1) begin
        trans_in_cnt_0 <= trans_in_cnt_0 + 16'h1;
    end
    else begin
        trans_in_cnt_0 <= trans_in_cnt_0;
    end
end

reg [15:0] trans_out_cnt_0;// for process Loop_VITIS_LOOP_67_1_proc39_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_0 <= 16'h0;
    end
    else if (Loop_VITIS_LOOP_67_1_proc39_U0.ap_done == 1'b1 && Loop_VITIS_LOOP_67_1_proc39_U0.ap_continue == 1'b1) begin
        trans_out_cnt_0 <= trans_out_cnt_0 + 16'h1;
    end
    else begin
        trans_out_cnt_0 <= trans_out_cnt_0;
    end
end

reg [15:0] trans_in_cnt_1;// for process myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_1 <= 16'h0;
    end
    else if (myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.start_write == 1'b1) begin
        trans_in_cnt_1 <= trans_in_cnt_1 + 16'h1;
    end
    else begin
        trans_in_cnt_1 <= trans_in_cnt_1;
    end
end

reg [15:0] trans_out_cnt_1;// for process myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_1 <= 16'h0;
    end
    else if (myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.ap_done == 1'b1 && myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.ap_continue == 1'b1) begin
        trans_out_cnt_1 <= trans_out_cnt_1 + 16'h1;
    end
    else begin
        trans_out_cnt_1 <= trans_out_cnt_1;
    end
end

reg [15:0] trans_in_cnt_2;// for process myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_2 <= 16'h0;
    end
    else if (myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.start_write == 1'b1) begin
        trans_in_cnt_2 <= trans_in_cnt_2 + 16'h1;
    end
    else begin
        trans_in_cnt_2 <= trans_in_cnt_2;
    end
end

reg [15:0] trans_out_cnt_2;// for process myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_2 <= 16'h0;
    end
    else if (myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.ap_done == 1'b1 && myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.ap_continue == 1'b1) begin
        trans_out_cnt_2 <= trans_out_cnt_2 + 16'h1;
    end
    else begin
        trans_out_cnt_2 <= trans_out_cnt_2;
    end
end

reg [15:0] trans_in_cnt_3;// for process myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_3 <= 16'h0;
    end
    else if (myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.start_write == 1'b1) begin
        trans_in_cnt_3 <= trans_in_cnt_3 + 16'h1;
    end
    else begin
        trans_in_cnt_3 <= trans_in_cnt_3;
    end
end

reg [15:0] trans_out_cnt_3;// for process myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_3 <= 16'h0;
    end
    else if (myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.ap_done == 1'b1 && myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.ap_continue == 1'b1) begin
        trans_out_cnt_3 <= trans_out_cnt_3 + 16'h1;
    end
    else begin
        trans_out_cnt_3 <= trans_out_cnt_3;
    end
end

reg [15:0] trans_in_cnt_4;// for process myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_4 <= 16'h0;
    end
    else if (myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.start_write == 1'b1) begin
        trans_in_cnt_4 <= trans_in_cnt_4 + 16'h1;
    end
    else begin
        trans_in_cnt_4 <= trans_in_cnt_4;
    end
end

reg [15:0] trans_out_cnt_4;// for process myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_4 <= 16'h0;
    end
    else if (myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.ap_done == 1'b1 && myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.ap_continue == 1'b1) begin
        trans_out_cnt_4 <= trans_out_cnt_4 + 16'h1;
    end
    else begin
        trans_out_cnt_4 <= trans_out_cnt_4;
    end
end

reg [15:0] trans_in_cnt_5;// for process myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_5 <= 16'h0;
    end
    else if (myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.start_write == 1'b1) begin
        trans_in_cnt_5 <= trans_in_cnt_5 + 16'h1;
    end
    else begin
        trans_in_cnt_5 <= trans_in_cnt_5;
    end
end

reg [15:0] trans_out_cnt_5;// for process myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_5 <= 16'h0;
    end
    else if (myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.ap_done == 1'b1 && myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.ap_continue == 1'b1) begin
        trans_out_cnt_5 <= trans_out_cnt_5 + 16'h1;
    end
    else begin
        trans_out_cnt_5 <= trans_out_cnt_5;
    end
end

reg [15:0] trans_in_cnt_6;// for process myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_6 <= 16'h0;
    end
    else if (myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.start_write == 1'b1) begin
        trans_in_cnt_6 <= trans_in_cnt_6 + 16'h1;
    end
    else begin
        trans_in_cnt_6 <= trans_in_cnt_6;
    end
end

reg [15:0] trans_out_cnt_6;// for process myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_6 <= 16'h0;
    end
    else if (myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.ap_done == 1'b1 && myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.ap_continue == 1'b1) begin
        trans_out_cnt_6 <= trans_out_cnt_6 + 16'h1;
    end
    else begin
        trans_out_cnt_6 <= trans_out_cnt_6;
    end
end

reg [15:0] trans_in_cnt_7;// for process myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_7 <= 16'h0;
    end
    else if (myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.start_write == 1'b1) begin
        trans_in_cnt_7 <= trans_in_cnt_7 + 16'h1;
    end
    else begin
        trans_in_cnt_7 <= trans_in_cnt_7;
    end
end

reg [15:0] trans_out_cnt_7;// for process myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_7 <= 16'h0;
    end
    else if (myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.ap_done == 1'b1 && myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.ap_continue == 1'b1) begin
        trans_out_cnt_7 <= trans_out_cnt_7 + 16'h1;
    end
    else begin
        trans_out_cnt_7 <= trans_out_cnt_7;
    end
end

reg [15:0] trans_in_cnt_8;// for process myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_8 <= 16'h0;
    end
    else if (myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.start_write == 1'b1) begin
        trans_in_cnt_8 <= trans_in_cnt_8 + 16'h1;
    end
    else begin
        trans_in_cnt_8 <= trans_in_cnt_8;
    end
end

reg [15:0] trans_out_cnt_8;// for process myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_8 <= 16'h0;
    end
    else if (myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.ap_done == 1'b1 && myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.ap_continue == 1'b1) begin
        trans_out_cnt_8 <= trans_out_cnt_8 + 16'h1;
    end
    else begin
        trans_out_cnt_8 <= trans_out_cnt_8;
    end
end

reg [15:0] trans_in_cnt_9;// for process myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_9 <= 16'h0;
    end
    else if (myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.start_write == 1'b1) begin
        trans_in_cnt_9 <= trans_in_cnt_9 + 16'h1;
    end
    else begin
        trans_in_cnt_9 <= trans_in_cnt_9;
    end
end

reg [15:0] trans_out_cnt_9;// for process myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_9 <= 16'h0;
    end
    else if (myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.ap_done == 1'b1 && myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.ap_continue == 1'b1) begin
        trans_out_cnt_9 <= trans_out_cnt_9 + 16'h1;
    end
    else begin
        trans_out_cnt_9 <= trans_out_cnt_9;
    end
end

reg [15:0] trans_in_cnt_10;// for process myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_10 <= 16'h0;
    end
    else if (myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.start_write == 1'b1) begin
        trans_in_cnt_10 <= trans_in_cnt_10 + 16'h1;
    end
    else begin
        trans_in_cnt_10 <= trans_in_cnt_10;
    end
end

reg [15:0] trans_out_cnt_10;// for process myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_10 <= 16'h0;
    end
    else if (myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.ap_done == 1'b1 && myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.ap_continue == 1'b1) begin
        trans_out_cnt_10 <= trans_out_cnt_10 + 16'h1;
    end
    else begin
        trans_out_cnt_10 <= trans_out_cnt_10;
    end
end

reg [15:0] trans_in_cnt_11;// for process myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_11 <= 16'h0;
    end
    else if (myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.start_write == 1'b1) begin
        trans_in_cnt_11 <= trans_in_cnt_11 + 16'h1;
    end
    else begin
        trans_in_cnt_11 <= trans_in_cnt_11;
    end
end

reg [15:0] trans_out_cnt_11;// for process myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_11 <= 16'h0;
    end
    else if (myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.ap_done == 1'b1 && myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.ap_continue == 1'b1) begin
        trans_out_cnt_11 <= trans_out_cnt_11 + 16'h1;
    end
    else begin
        trans_out_cnt_11 <= trans_out_cnt_11;
    end
end

reg [15:0] trans_in_cnt_12;// for process myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_12 <= 16'h0;
    end
    else if (myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.start_write == 1'b1) begin
        trans_in_cnt_12 <= trans_in_cnt_12 + 16'h1;
    end
    else begin
        trans_in_cnt_12 <= trans_in_cnt_12;
    end
end

reg [15:0] trans_out_cnt_12;// for process myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_12 <= 16'h0;
    end
    else if (myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.ap_done == 1'b1 && myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.ap_continue == 1'b1) begin
        trans_out_cnt_12 <= trans_out_cnt_12 + 16'h1;
    end
    else begin
        trans_out_cnt_12 <= trans_out_cnt_12;
    end
end

reg [15:0] trans_in_cnt_13;// for process myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_13 <= 16'h0;
    end
    else if (myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.start_write == 1'b1) begin
        trans_in_cnt_13 <= trans_in_cnt_13 + 16'h1;
    end
    else begin
        trans_in_cnt_13 <= trans_in_cnt_13;
    end
end

reg [15:0] trans_out_cnt_13;// for process myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_13 <= 16'h0;
    end
    else if (myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.ap_done == 1'b1 && myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.ap_continue == 1'b1) begin
        trans_out_cnt_13 <= trans_out_cnt_13 + 16'h1;
    end
    else begin
        trans_out_cnt_13 <= trans_out_cnt_13;
    end
end

reg [15:0] trans_in_cnt_14;// for process myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_14 <= 16'h0;
    end
    else if (myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.start_write == 1'b1) begin
        trans_in_cnt_14 <= trans_in_cnt_14 + 16'h1;
    end
    else begin
        trans_in_cnt_14 <= trans_in_cnt_14;
    end
end

reg [15:0] trans_out_cnt_14;// for process myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_14 <= 16'h0;
    end
    else if (myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.ap_done == 1'b1 && myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.ap_continue == 1'b1) begin
        trans_out_cnt_14 <= trans_out_cnt_14 + 16'h1;
    end
    else begin
        trans_out_cnt_14 <= trans_out_cnt_14;
    end
end

reg [15:0] trans_in_cnt_15;// for process myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_15 <= 16'h0;
    end
    else if (myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.start_write == 1'b1) begin
        trans_in_cnt_15 <= trans_in_cnt_15 + 16'h1;
    end
    else begin
        trans_in_cnt_15 <= trans_in_cnt_15;
    end
end

reg [15:0] trans_out_cnt_15;// for process myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_15 <= 16'h0;
    end
    else if (myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.ap_done == 1'b1 && myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.ap_continue == 1'b1) begin
        trans_out_cnt_15 <= trans_out_cnt_15 + 16'h1;
    end
    else begin
        trans_out_cnt_15 <= trans_out_cnt_15;
    end
end

reg [15:0] trans_in_cnt_16;// for process myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_16 <= 16'h0;
    end
    else if (myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.start_write == 1'b1) begin
        trans_in_cnt_16 <= trans_in_cnt_16 + 16'h1;
    end
    else begin
        trans_in_cnt_16 <= trans_in_cnt_16;
    end
end

reg [15:0] trans_out_cnt_16;// for process myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_16 <= 16'h0;
    end
    else if (myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.ap_done == 1'b1 && myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.ap_continue == 1'b1) begin
        trans_out_cnt_16 <= trans_out_cnt_16 + 16'h1;
    end
    else begin
        trans_out_cnt_16 <= trans_out_cnt_16;
    end
end

reg [15:0] trans_in_cnt_17;// for process myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_17 <= 16'h0;
    end
    else if (myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.start_write == 1'b1) begin
        trans_in_cnt_17 <= trans_in_cnt_17 + 16'h1;
    end
    else begin
        trans_in_cnt_17 <= trans_in_cnt_17;
    end
end

reg [15:0] trans_out_cnt_17;// for process myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_17 <= 16'h0;
    end
    else if (myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.ap_done == 1'b1 && myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.ap_continue == 1'b1) begin
        trans_out_cnt_17 <= trans_out_cnt_17 + 16'h1;
    end
    else begin
        trans_out_cnt_17 <= trans_out_cnt_17;
    end
end

reg [15:0] trans_in_cnt_18;// for process myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config23_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_18 <= 16'h0;
    end
    else if (myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config23_U0.start_write == 1'b1) begin
        trans_in_cnt_18 <= trans_in_cnt_18 + 16'h1;
    end
    else begin
        trans_in_cnt_18 <= trans_in_cnt_18;
    end
end

reg [15:0] trans_out_cnt_18;// for process myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config23_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_18 <= 16'h0;
    end
    else if (myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config23_U0.ap_done == 1'b1 && myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config23_U0.ap_continue == 1'b1) begin
        trans_out_cnt_18 <= trans_out_cnt_18 + 16'h1;
    end
    else begin
        trans_out_cnt_18 <= trans_out_cnt_18;
    end
end

reg [15:0] trans_in_cnt_19;// for process entry_proc_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_19 <= 16'h0;
    end
    else if (entry_proc_U0.start_write == 1'b1) begin
        trans_in_cnt_19 <= trans_in_cnt_19 + 16'h1;
    end
    else begin
        trans_in_cnt_19 <= trans_in_cnt_19;
    end
end

reg [15:0] trans_out_cnt_19;// for process entry_proc_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_19 <= 16'h0;
    end
    else if (entry_proc_U0.ap_done == 1'b1 && entry_proc_U0.ap_continue == 1'b1) begin
        trans_out_cnt_19 <= trans_out_cnt_19 + 16'h1;
    end
    else begin
        trans_out_cnt_19 <= trans_out_cnt_19;
    end
end

    // Process: entry_proc_U0
    alveo_hls4ml_hls_deadlock_detect_unit #(26, 0, 3, 3) alveo_hls4ml_hls_deadlock_detect_unit_0 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_0),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_0),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_0),
        .token_in_vec(token_in_vec_0),
        .dl_detect_in(dl_detect_out),
        .origin(origin[0]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_0),
        .out_chan_dep_data(out_chan_dep_data_0),
        .token_out_vec(token_out_vec_0),
        .dl_detect_out(dl_in_vec[0]));

    assign proc_0_data_FIFO_blk[0] = 1'b0 | (~entry_proc_U0.out_r_c_blk_n);
    assign proc_0_data_PIPO_blk[0] = 1'b0;
    assign proc_0_start_FIFO_blk[0] = 1'b0 | (~start_for_Loop_VITIS_LOOP_93_5_proc41_U0_U.if_full_n & entry_proc_U0.ap_start & ~entry_proc_U0.real_start & (trans_in_cnt_19 == trans_out_cnt_19) & ~start_for_Loop_VITIS_LOOP_93_5_proc41_U0_U.if_read);
    assign proc_0_TLF_FIFO_blk[0] = 1'b0;
    assign proc_0_input_sync_blk[0] = 1'b0;
    assign proc_0_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_0[0] = dl_detect_out ? proc_dep_vld_vec_0_reg[0] : (proc_0_data_FIFO_blk[0] | proc_0_data_PIPO_blk[0] | proc_0_start_FIFO_blk[0] | proc_0_TLF_FIFO_blk[0] | proc_0_input_sync_blk[0] | proc_0_output_sync_blk[0]);
    assign proc_0_data_FIFO_blk[1] = 1'b0;
    assign proc_0_data_PIPO_blk[1] = 1'b0;
    assign proc_0_start_FIFO_blk[1] = 1'b0;
    assign proc_0_TLF_FIFO_blk[1] = 1'b0;
    assign proc_0_input_sync_blk[1] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_Loop_VITIS_LOOP_67_1_proc39_U0_ap_ready);
    assign proc_0_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_0[1] = dl_detect_out ? proc_dep_vld_vec_0_reg[1] : (proc_0_data_FIFO_blk[1] | proc_0_data_PIPO_blk[1] | proc_0_start_FIFO_blk[1] | proc_0_TLF_FIFO_blk[1] | proc_0_input_sync_blk[1] | proc_0_output_sync_blk[1]);
    assign proc_0_data_FIFO_blk[2] = 1'b0;
    assign proc_0_data_PIPO_blk[2] = 1'b0;
    assign proc_0_start_FIFO_blk[2] = 1'b0;
    assign proc_0_TLF_FIFO_blk[2] = 1'b0;
    assign proc_0_input_sync_blk[2] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_Loop_VITIS_LOOP_74_3_proc40_U0_ap_ready);
    assign proc_0_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_0[2] = dl_detect_out ? proc_dep_vld_vec_0_reg[2] : (proc_0_data_FIFO_blk[2] | proc_0_data_PIPO_blk[2] | proc_0_start_FIFO_blk[2] | proc_0_TLF_FIFO_blk[2] | proc_0_input_sync_blk[2] | proc_0_output_sync_blk[2]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_0_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_0_reg <= proc_dep_vld_vec_0;
        end
    end
    assign in_chan_dep_vld_vec_0[0] = dep_chan_vld_1_0;
    assign in_chan_dep_data_vec_0[25 : 0] = dep_chan_data_1_0;
    assign token_in_vec_0[0] = token_1_0;
    assign in_chan_dep_vld_vec_0[1] = dep_chan_vld_2_0;
    assign in_chan_dep_data_vec_0[51 : 26] = dep_chan_data_2_0;
    assign token_in_vec_0[1] = token_2_0;
    assign in_chan_dep_vld_vec_0[2] = dep_chan_vld_25_0;
    assign in_chan_dep_data_vec_0[77 : 52] = dep_chan_data_25_0;
    assign token_in_vec_0[2] = token_25_0;
    assign dep_chan_vld_0_25 = out_chan_dep_vld_vec_0[0];
    assign dep_chan_data_0_25 = out_chan_dep_data_0;
    assign token_0_25 = token_out_vec_0[0];
    assign dep_chan_vld_0_1 = out_chan_dep_vld_vec_0[1];
    assign dep_chan_data_0_1 = out_chan_dep_data_0;
    assign token_0_1 = token_out_vec_0[1];
    assign dep_chan_vld_0_2 = out_chan_dep_vld_vec_0[2];
    assign dep_chan_data_0_2 = out_chan_dep_data_0;
    assign token_0_2 = token_out_vec_0[2];

    // Process: Loop_VITIS_LOOP_67_1_proc39_U0
    alveo_hls4ml_hls_deadlock_detect_unit #(26, 1, 4, 4) alveo_hls4ml_hls_deadlock_detect_unit_1 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_1),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_1),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_1),
        .token_in_vec(token_in_vec_1),
        .dl_detect_in(dl_detect_out),
        .origin(origin[1]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_1),
        .out_chan_dep_data(out_chan_dep_data_1),
        .token_out_vec(token_out_vec_1),
        .dl_detect_out(dl_in_vec[1]));

    assign proc_1_data_FIFO_blk[0] = 1'b0 | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_0_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_1_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_2_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_3_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_4_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_5_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_6_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_7_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_8_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_9_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_10_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_11_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_12_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_13_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_14_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_15_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_16_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_17_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_18_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_19_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_20_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_21_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_22_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_23_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_24_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_25_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_26_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_27_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_28_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_29_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_30_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_31_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_32_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_33_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_34_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_35_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_36_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_37_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_38_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_39_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_40_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_41_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_42_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_43_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_44_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_45_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_46_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_47_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_48_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_49_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_50_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_51_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_52_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_53_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_54_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_55_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_56_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_57_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_58_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_59_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_60_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_61_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_62_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_63_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_64_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_65_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_66_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_67_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_68_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_69_blk_n);
    assign proc_1_data_PIPO_blk[0] = 1'b0;
    assign proc_1_start_FIFO_blk[0] = 1'b0 | (~start_for_myproject_U0_U.if_full_n & Loop_VITIS_LOOP_67_1_proc39_U0.ap_start & ~Loop_VITIS_LOOP_67_1_proc39_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_myproject_U0_U.if_read);
    assign proc_1_TLF_FIFO_blk[0] = 1'b0;
    assign proc_1_input_sync_blk[0] = 1'b0;
    assign proc_1_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_1[0] = dl_detect_out ? proc_dep_vld_vec_1_reg[0] : (proc_1_data_FIFO_blk[0] | proc_1_data_PIPO_blk[0] | proc_1_start_FIFO_blk[0] | proc_1_TLF_FIFO_blk[0] | proc_1_input_sync_blk[0] | proc_1_output_sync_blk[0]);
    assign proc_1_data_FIFO_blk[1] = 1'b0 | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_0_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_1_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_2_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_3_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_4_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_5_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_6_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_7_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_8_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_9_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_10_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_11_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_12_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_13_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_14_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_15_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_16_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_17_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_18_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_19_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_20_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_21_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_22_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_23_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_24_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_25_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_26_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_27_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_28_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_29_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_30_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_31_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_32_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_33_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_34_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_35_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_36_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_37_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_38_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_39_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_40_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_41_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_42_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_43_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_44_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_45_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_46_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_47_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_48_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_49_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_50_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_51_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_52_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_53_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_54_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_55_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_56_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_57_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_58_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_59_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_60_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_61_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_62_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_63_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_64_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_65_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_66_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_67_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_68_blk_n) | (~Loop_VITIS_LOOP_67_1_proc39_U0.grp_Loop_VITIS_LOOP_67_1_proc39_Pipeline_VITIS_LOOP_67_1_VITIS_LOOP_68_2_fu_193.in_stream1_69_blk_n);
    assign proc_1_data_PIPO_blk[1] = 1'b0;
    assign proc_1_start_FIFO_blk[1] = 1'b0;
    assign proc_1_TLF_FIFO_blk[1] = 1'b0;
    assign proc_1_input_sync_blk[1] = 1'b0;
    assign proc_1_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_1[1] = dl_detect_out ? proc_dep_vld_vec_1_reg[1] : (proc_1_data_FIFO_blk[1] | proc_1_data_PIPO_blk[1] | proc_1_start_FIFO_blk[1] | proc_1_TLF_FIFO_blk[1] | proc_1_input_sync_blk[1] | proc_1_output_sync_blk[1]);
    assign proc_1_data_FIFO_blk[2] = 1'b0;
    assign proc_1_data_PIPO_blk[2] = 1'b0;
    assign proc_1_start_FIFO_blk[2] = 1'b0;
    assign proc_1_TLF_FIFO_blk[2] = 1'b0;
    assign proc_1_input_sync_blk[2] = 1'b0 | (ap_sync_Loop_VITIS_LOOP_67_1_proc39_U0_ap_ready & Loop_VITIS_LOOP_67_1_proc39_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_1_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_1[2] = dl_detect_out ? proc_dep_vld_vec_1_reg[2] : (proc_1_data_FIFO_blk[2] | proc_1_data_PIPO_blk[2] | proc_1_start_FIFO_blk[2] | proc_1_TLF_FIFO_blk[2] | proc_1_input_sync_blk[2] | proc_1_output_sync_blk[2]);
    assign proc_1_data_FIFO_blk[3] = 1'b0;
    assign proc_1_data_PIPO_blk[3] = 1'b0;
    assign proc_1_start_FIFO_blk[3] = 1'b0;
    assign proc_1_TLF_FIFO_blk[3] = 1'b0;
    assign proc_1_input_sync_blk[3] = 1'b0 | (ap_sync_Loop_VITIS_LOOP_67_1_proc39_U0_ap_ready & Loop_VITIS_LOOP_67_1_proc39_U0.ap_idle & ~ap_sync_Loop_VITIS_LOOP_74_3_proc40_U0_ap_ready);
    assign proc_1_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_1[3] = dl_detect_out ? proc_dep_vld_vec_1_reg[3] : (proc_1_data_FIFO_blk[3] | proc_1_data_PIPO_blk[3] | proc_1_start_FIFO_blk[3] | proc_1_TLF_FIFO_blk[3] | proc_1_input_sync_blk[3] | proc_1_output_sync_blk[3]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_1_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_1_reg <= proc_dep_vld_vec_1;
        end
    end
    assign in_chan_dep_vld_vec_1[0] = dep_chan_vld_0_1;
    assign in_chan_dep_data_vec_1[25 : 0] = dep_chan_data_0_1;
    assign token_in_vec_1[0] = token_0_1;
    assign in_chan_dep_vld_vec_1[1] = dep_chan_vld_2_1;
    assign in_chan_dep_data_vec_1[51 : 26] = dep_chan_data_2_1;
    assign token_in_vec_1[1] = token_2_1;
    assign in_chan_dep_vld_vec_1[2] = dep_chan_vld_3_1;
    assign in_chan_dep_data_vec_1[77 : 52] = dep_chan_data_3_1;
    assign token_in_vec_1[2] = token_3_1;
    assign in_chan_dep_vld_vec_1[3] = dep_chan_vld_4_1;
    assign in_chan_dep_data_vec_1[103 : 78] = dep_chan_data_4_1;
    assign token_in_vec_1[3] = token_4_1;
    assign dep_chan_vld_1_3 = out_chan_dep_vld_vec_1[0];
    assign dep_chan_data_1_3 = out_chan_dep_data_1;
    assign token_1_3 = token_out_vec_1[0];
    assign dep_chan_vld_1_4 = out_chan_dep_vld_vec_1[1];
    assign dep_chan_data_1_4 = out_chan_dep_data_1;
    assign token_1_4 = token_out_vec_1[1];
    assign dep_chan_vld_1_0 = out_chan_dep_vld_vec_1[2];
    assign dep_chan_data_1_0 = out_chan_dep_data_1;
    assign token_1_0 = token_out_vec_1[2];
    assign dep_chan_vld_1_2 = out_chan_dep_vld_vec_1[3];
    assign dep_chan_data_1_2 = out_chan_dep_data_1;
    assign token_1_2 = token_out_vec_1[3];

    // Process: Loop_VITIS_LOOP_74_3_proc40_U0
    alveo_hls4ml_hls_deadlock_detect_unit #(26, 2, 4, 4) alveo_hls4ml_hls_deadlock_detect_unit_2 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_2),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_2),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_2),
        .token_in_vec(token_in_vec_2),
        .dl_detect_in(dl_detect_out),
        .origin(origin[2]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_2),
        .out_chan_dep_data(out_chan_dep_data_2),
        .token_out_vec(token_out_vec_2),
        .dl_detect_out(dl_in_vec[2]));

    assign proc_2_data_FIFO_blk[0] = 1'b0 | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_0_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_1_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_2_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_3_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_4_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_5_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_6_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_7_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_8_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_9_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_10_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_11_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_12_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_13_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_14_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_15_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_16_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_17_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_18_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_19_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_20_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_21_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_22_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_23_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_24_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_25_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_26_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_27_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_28_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_29_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_30_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_31_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_32_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_33_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_34_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_35_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_36_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_37_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_38_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_39_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_40_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_41_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_42_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_43_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_44_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_45_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_46_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_47_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_48_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_49_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_50_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_51_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_52_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_53_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_54_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_55_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_56_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_57_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_58_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_59_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_60_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_61_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_62_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_63_blk_n);
    assign proc_2_data_PIPO_blk[0] = 1'b0;
    assign proc_2_start_FIFO_blk[0] = 1'b0;
    assign proc_2_TLF_FIFO_blk[0] = 1'b0;
    assign proc_2_input_sync_blk[0] = 1'b0;
    assign proc_2_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_2[0] = dl_detect_out ? proc_dep_vld_vec_2_reg[0] : (proc_2_data_FIFO_blk[0] | proc_2_data_PIPO_blk[0] | proc_2_start_FIFO_blk[0] | proc_2_TLF_FIFO_blk[0] | proc_2_input_sync_blk[0] | proc_2_output_sync_blk[0]);
    assign proc_2_data_FIFO_blk[1] = 1'b0 | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_0_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_1_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_2_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_3_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_4_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_5_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_6_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_7_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_8_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_9_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_10_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_11_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_12_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_13_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_14_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_15_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_16_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_17_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_18_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_19_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_20_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_21_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_22_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_23_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_24_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_25_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_26_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_27_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_28_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_29_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_30_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_31_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_32_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_33_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_34_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_35_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_36_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_37_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_38_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_39_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_40_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_41_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_42_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_43_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_44_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_45_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_46_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_47_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_48_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_49_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_50_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_51_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_52_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_53_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_54_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_55_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_56_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_57_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_58_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_59_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_60_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_61_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_62_blk_n) | (~Loop_VITIS_LOOP_74_3_proc40_U0.grp_Loop_VITIS_LOOP_74_3_proc40_Pipeline_VITIS_LOOP_74_3_VITIS_LOOP_75_4_fu_181.in_stream2_63_blk_n);
    assign proc_2_data_PIPO_blk[1] = 1'b0;
    assign proc_2_start_FIFO_blk[1] = 1'b0;
    assign proc_2_TLF_FIFO_blk[1] = 1'b0;
    assign proc_2_input_sync_blk[1] = 1'b0;
    assign proc_2_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_2[1] = dl_detect_out ? proc_dep_vld_vec_2_reg[1] : (proc_2_data_FIFO_blk[1] | proc_2_data_PIPO_blk[1] | proc_2_start_FIFO_blk[1] | proc_2_TLF_FIFO_blk[1] | proc_2_input_sync_blk[1] | proc_2_output_sync_blk[1]);
    assign proc_2_data_FIFO_blk[2] = 1'b0;
    assign proc_2_data_PIPO_blk[2] = 1'b0;
    assign proc_2_start_FIFO_blk[2] = 1'b0;
    assign proc_2_TLF_FIFO_blk[2] = 1'b0;
    assign proc_2_input_sync_blk[2] = 1'b0 | (ap_sync_Loop_VITIS_LOOP_74_3_proc40_U0_ap_ready & Loop_VITIS_LOOP_74_3_proc40_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_2_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_2[2] = dl_detect_out ? proc_dep_vld_vec_2_reg[2] : (proc_2_data_FIFO_blk[2] | proc_2_data_PIPO_blk[2] | proc_2_start_FIFO_blk[2] | proc_2_TLF_FIFO_blk[2] | proc_2_input_sync_blk[2] | proc_2_output_sync_blk[2]);
    assign proc_2_data_FIFO_blk[3] = 1'b0;
    assign proc_2_data_PIPO_blk[3] = 1'b0;
    assign proc_2_start_FIFO_blk[3] = 1'b0;
    assign proc_2_TLF_FIFO_blk[3] = 1'b0;
    assign proc_2_input_sync_blk[3] = 1'b0 | (ap_sync_Loop_VITIS_LOOP_74_3_proc40_U0_ap_ready & Loop_VITIS_LOOP_74_3_proc40_U0.ap_idle & ~ap_sync_Loop_VITIS_LOOP_67_1_proc39_U0_ap_ready);
    assign proc_2_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_2[3] = dl_detect_out ? proc_dep_vld_vec_2_reg[3] : (proc_2_data_FIFO_blk[3] | proc_2_data_PIPO_blk[3] | proc_2_start_FIFO_blk[3] | proc_2_TLF_FIFO_blk[3] | proc_2_input_sync_blk[3] | proc_2_output_sync_blk[3]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_2_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_2_reg <= proc_dep_vld_vec_2;
        end
    end
    assign in_chan_dep_vld_vec_2[0] = dep_chan_vld_0_2;
    assign in_chan_dep_data_vec_2[25 : 0] = dep_chan_data_0_2;
    assign token_in_vec_2[0] = token_0_2;
    assign in_chan_dep_vld_vec_2[1] = dep_chan_vld_1_2;
    assign in_chan_dep_data_vec_2[51 : 26] = dep_chan_data_1_2;
    assign token_in_vec_2[1] = token_1_2;
    assign in_chan_dep_vld_vec_2[2] = dep_chan_vld_3_2;
    assign in_chan_dep_data_vec_2[77 : 52] = dep_chan_data_3_2;
    assign token_in_vec_2[2] = token_3_2;
    assign in_chan_dep_vld_vec_2[3] = dep_chan_vld_20_2;
    assign in_chan_dep_data_vec_2[103 : 78] = dep_chan_data_20_2;
    assign token_in_vec_2[3] = token_20_2;
    assign dep_chan_vld_2_3 = out_chan_dep_vld_vec_2[0];
    assign dep_chan_data_2_3 = out_chan_dep_data_2;
    assign token_2_3 = token_out_vec_2[0];
    assign dep_chan_vld_2_20 = out_chan_dep_vld_vec_2[1];
    assign dep_chan_data_2_20 = out_chan_dep_data_2;
    assign token_2_20 = token_out_vec_2[1];
    assign dep_chan_vld_2_0 = out_chan_dep_vld_vec_2[2];
    assign dep_chan_data_2_0 = out_chan_dep_data_2;
    assign token_2_0 = token_out_vec_2[2];
    assign dep_chan_vld_2_1 = out_chan_dep_vld_vec_2[3];
    assign dep_chan_data_2_1 = out_chan_dep_data_2;
    assign token_2_1 = token_out_vec_2[3];

    // Process: myproject_U0
    alveo_hls4ml_hls_deadlock_detect_unit #(26, 3, 3, 3) alveo_hls4ml_hls_deadlock_detect_unit_3 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_3),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_3),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_3),
        .token_in_vec(token_in_vec_3),
        .dl_detect_in(dl_detect_out),
        .origin(origin[3]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_3),
        .out_chan_dep_data(out_chan_dep_data_3),
        .token_out_vec(token_out_vec_3),
        .dl_detect_out(dl_in_vec[3]));

    assign proc_3_data_FIFO_blk[0] = 1'b0 | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_0_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_1_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_2_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_3_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_4_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_5_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_6_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_7_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_8_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_9_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_10_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_11_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_12_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_13_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_14_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_15_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_16_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_17_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_18_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_19_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_20_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_21_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_22_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_23_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_24_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_25_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_26_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_27_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_28_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_29_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_30_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_31_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_32_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_33_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_34_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_35_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_36_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_37_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_38_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_39_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_40_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_41_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_42_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_43_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_44_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_45_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_46_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_47_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_48_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_49_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_50_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_51_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_52_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_53_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_54_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_55_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_56_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_57_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_58_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_59_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_60_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_61_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_62_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_63_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_64_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_65_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_66_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_67_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_68_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_69_blk_n);
    assign proc_3_data_PIPO_blk[0] = 1'b0;
    assign proc_3_start_FIFO_blk[0] = 1'b0 | (~start_for_myproject_U0_U.if_empty_n & myproject_U0.ap_idle & ~start_for_myproject_U0_U.if_write);
    assign proc_3_TLF_FIFO_blk[0] = 1'b0;
    assign proc_3_input_sync_blk[0] = 1'b0;
    assign proc_3_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_3[0] = dl_detect_out ? proc_dep_vld_vec_3_reg[0] : (proc_3_data_FIFO_blk[0] | proc_3_data_PIPO_blk[0] | proc_3_start_FIFO_blk[0] | proc_3_TLF_FIFO_blk[0] | proc_3_input_sync_blk[0] | proc_3_output_sync_blk[0]);
    assign proc_3_data_FIFO_blk[1] = 1'b0 | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_0_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_1_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_2_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_3_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_4_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_5_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_6_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_7_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_8_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_9_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_10_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_11_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_12_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_13_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_14_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_15_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_16_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_17_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_18_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_19_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_20_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_21_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_22_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_23_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_24_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_25_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_26_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_27_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_28_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_29_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_30_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_31_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_32_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_33_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_34_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_35_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_36_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_37_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_38_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_39_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_40_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_41_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_42_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_43_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_44_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_45_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_46_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_47_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_48_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_49_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_50_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_51_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_52_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_53_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_54_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_55_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_56_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_57_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_58_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_59_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_60_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_61_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_62_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_63_blk_n);
    assign proc_3_data_PIPO_blk[1] = 1'b0;
    assign proc_3_start_FIFO_blk[1] = 1'b0;
    assign proc_3_TLF_FIFO_blk[1] = 1'b0;
    assign proc_3_input_sync_blk[1] = 1'b0;
    assign proc_3_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_3[1] = dl_detect_out ? proc_dep_vld_vec_3_reg[1] : (proc_3_data_FIFO_blk[1] | proc_3_data_PIPO_blk[1] | proc_3_start_FIFO_blk[1] | proc_3_TLF_FIFO_blk[1] | proc_3_input_sync_blk[1] | proc_3_output_sync_blk[1]);
    assign proc_3_data_FIFO_blk[2] = 1'b0 | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_0_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_1_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_2_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_3_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_4_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_5_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_6_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_7_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_8_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_9_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_10_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_11_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_12_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_13_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_14_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_15_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_16_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_17_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_18_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_19_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_20_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_21_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_22_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_23_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_24_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_25_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_26_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_27_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_28_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_29_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_30_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_31_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_32_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_33_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_34_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_35_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_36_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_37_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_38_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_39_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_40_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_41_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_42_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_43_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_44_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_45_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_46_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_47_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_48_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_49_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_50_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_51_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_52_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_53_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_54_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_55_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_56_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_57_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_58_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_59_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_60_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_61_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_62_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_63_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_64_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_65_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_66_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_67_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_68_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_69_blk_n);
    assign proc_3_data_PIPO_blk[2] = 1'b0;
    assign proc_3_start_FIFO_blk[2] = 1'b0;
    assign proc_3_TLF_FIFO_blk[2] = 1'b0;
    assign proc_3_input_sync_blk[2] = 1'b0;
    assign proc_3_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_3[2] = dl_detect_out ? proc_dep_vld_vec_3_reg[2] : (proc_3_data_FIFO_blk[2] | proc_3_data_PIPO_blk[2] | proc_3_start_FIFO_blk[2] | proc_3_TLF_FIFO_blk[2] | proc_3_input_sync_blk[2] | proc_3_output_sync_blk[2]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_3_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_3_reg <= proc_dep_vld_vec_3;
        end
    end
    assign in_chan_dep_vld_vec_3[0] = dep_chan_vld_1_3;
    assign in_chan_dep_data_vec_3[25 : 0] = dep_chan_data_1_3;
    assign token_in_vec_3[0] = token_1_3;
    assign in_chan_dep_vld_vec_3[1] = dep_chan_vld_2_3;
    assign in_chan_dep_data_vec_3[51 : 26] = dep_chan_data_2_3;
    assign token_in_vec_3[1] = token_2_3;
    assign in_chan_dep_vld_vec_3[2] = dep_chan_vld_25_3;
    assign in_chan_dep_data_vec_3[77 : 52] = dep_chan_data_25_3;
    assign token_in_vec_3[2] = token_25_3;
    assign dep_chan_vld_3_1 = out_chan_dep_vld_vec_3[0];
    assign dep_chan_data_3_1 = out_chan_dep_data_3;
    assign token_3_1 = token_out_vec_3[0];
    assign dep_chan_vld_3_2 = out_chan_dep_vld_vec_3[1];
    assign dep_chan_data_3_2 = out_chan_dep_data_3;
    assign token_3_2 = token_out_vec_3[1];
    assign dep_chan_vld_3_25 = out_chan_dep_vld_vec_3[2];
    assign dep_chan_data_3_25 = out_chan_dep_data_3;
    assign token_3_25 = token_out_vec_3[2];

    // Process: myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0
    alveo_hls4ml_hls_deadlock_detect_unit #(26, 4, 2, 2) alveo_hls4ml_hls_deadlock_detect_unit_4 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_4),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_4),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_4),
        .token_in_vec(token_in_vec_4),
        .dl_detect_in(dl_detect_out),
        .origin(origin[4]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_4),
        .out_chan_dep_data(out_chan_dep_data_4),
        .token_out_vec(token_out_vec_4),
        .dl_detect_out(dl_in_vec[4]));

    assign proc_4_data_FIFO_blk[0] = 1'b0 | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_0_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_1_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_2_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_3_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_4_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_5_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_6_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_7_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_8_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_9_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_10_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_11_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_12_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_13_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_14_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_15_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_16_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_17_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_18_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_19_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_20_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_21_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_22_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_23_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_24_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_25_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_26_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_27_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_28_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_29_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_30_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_31_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_32_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_33_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_34_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_35_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_36_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_37_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_38_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_39_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_40_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_41_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_42_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_43_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_44_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_45_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_46_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_47_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_48_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_49_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_50_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_51_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_52_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_53_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_54_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_55_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_56_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_57_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_58_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_59_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_60_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_61_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_62_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_63_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_64_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_65_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_66_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_67_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_68_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.grp_bidirectional_array_ap_fixed_ap_fixed_config2_Pipeline_VITIS_LOOP_111_1_fu_2138.in_stream1_69_blk_n);
    assign proc_4_data_PIPO_blk[0] = 1'b0;
    assign proc_4_start_FIFO_blk[0] = 1'b0;
    assign proc_4_TLF_FIFO_blk[0] = 1'b0;
    assign proc_4_input_sync_blk[0] = 1'b0;
    assign proc_4_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_4[0] = dl_detect_out ? proc_dep_vld_vec_4_reg[0] : (proc_4_data_FIFO_blk[0] | proc_4_data_PIPO_blk[0] | proc_4_start_FIFO_blk[0] | proc_4_TLF_FIFO_blk[0] | proc_4_input_sync_blk[0] | proc_4_output_sync_blk[0]);
    assign proc_4_data_FIFO_blk[1] = 1'b0 | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_0_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_1_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_2_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_3_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_4_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_5_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_6_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_7_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_8_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_9_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_10_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_11_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_12_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_13_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_14_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_15_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_16_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_17_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_18_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_19_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_20_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_21_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_22_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_23_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_24_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_25_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_26_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_27_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_28_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_29_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_30_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_31_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_32_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_33_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_34_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_35_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_36_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_37_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_38_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_39_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_40_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_41_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_42_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_43_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_44_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_45_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_46_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_47_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_48_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_49_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_50_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_51_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_52_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_53_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_54_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_55_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_56_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_57_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_58_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_59_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_60_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_61_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_62_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_63_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_64_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_65_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_66_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_67_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_68_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_69_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_70_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_71_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_72_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_73_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_74_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_75_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_76_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_77_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_78_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_79_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_80_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_81_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_82_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_83_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_84_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_85_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_86_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_87_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_88_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_89_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_90_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_91_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_92_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_93_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_94_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_95_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_96_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_97_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_98_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_99_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_100_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_101_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_102_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_103_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_104_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_105_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_106_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_107_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_108_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_109_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_110_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_111_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_112_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_113_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_114_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_115_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_116_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_117_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_118_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_119_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_120_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_121_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_122_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_123_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_124_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_125_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_126_blk_n) | (~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.layer2_out_127_blk_n);
    assign proc_4_data_PIPO_blk[1] = 1'b0;
    assign proc_4_start_FIFO_blk[1] = 1'b0 | (~myproject_U0.start_for_linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0_U.if_full_n & myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.ap_start & ~myproject_U0.bidirectional_array_ap_fixed_16_6_5_3_0_ap_fixed_33_4_5_3_0_config2_U0.real_start & (trans_in_cnt_1 == trans_out_cnt_1) & ~myproject_U0.start_for_linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0_U.if_read);
    assign proc_4_TLF_FIFO_blk[1] = 1'b0;
    assign proc_4_input_sync_blk[1] = 1'b0;
    assign proc_4_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_4[1] = dl_detect_out ? proc_dep_vld_vec_4_reg[1] : (proc_4_data_FIFO_blk[1] | proc_4_data_PIPO_blk[1] | proc_4_start_FIFO_blk[1] | proc_4_TLF_FIFO_blk[1] | proc_4_input_sync_blk[1] | proc_4_output_sync_blk[1]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_4_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_4_reg <= proc_dep_vld_vec_4;
        end
    end
    assign in_chan_dep_vld_vec_4[0] = dep_chan_vld_1_4;
    assign in_chan_dep_data_vec_4[25 : 0] = dep_chan_data_1_4;
    assign token_in_vec_4[0] = token_1_4;
    assign in_chan_dep_vld_vec_4[1] = dep_chan_vld_5_4;
    assign in_chan_dep_data_vec_4[51 : 26] = dep_chan_data_5_4;
    assign token_in_vec_4[1] = token_5_4;
    assign dep_chan_vld_4_1 = out_chan_dep_vld_vec_4[0];
    assign dep_chan_data_4_1 = out_chan_dep_data_4;
    assign token_4_1 = token_out_vec_4[0];
    assign dep_chan_vld_4_5 = out_chan_dep_vld_vec_4[1];
    assign dep_chan_data_4_5 = out_chan_dep_data_4;
    assign token_4_5 = token_out_vec_4[1];

    // Process: myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0
    alveo_hls4ml_hls_deadlock_detect_unit #(26, 5, 2, 2) alveo_hls4ml_hls_deadlock_detect_unit_5 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_5),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_5),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_5),
        .token_in_vec(token_in_vec_5),
        .dl_detect_in(dl_detect_out),
        .origin(origin[5]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_5),
        .out_chan_dep_data(out_chan_dep_data_5),
        .token_out_vec(token_out_vec_5),
        .dl_detect_out(dl_in_vec[5]));

    assign proc_5_data_FIFO_blk[0] = 1'b0 | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_0_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_1_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_2_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_3_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_4_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_5_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_6_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_7_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_8_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_9_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_10_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_11_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_12_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_13_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_14_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_15_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_16_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_17_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_18_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_19_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_20_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_21_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_22_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_23_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_24_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_25_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_26_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_27_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_28_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_29_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_30_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_31_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_32_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_33_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_34_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_35_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_36_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_37_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_38_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_39_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_40_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_41_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_42_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_43_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_44_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_45_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_46_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_47_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_48_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_49_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_50_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_51_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_52_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_53_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_54_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_55_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_56_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_57_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_58_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_59_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_60_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_61_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_62_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_63_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_64_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_65_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_66_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_67_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_68_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_69_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_70_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_71_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_72_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_73_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_74_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_75_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_76_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_77_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_78_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_79_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_80_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_81_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_82_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_83_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_84_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_85_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_86_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_87_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_88_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_89_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_90_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_91_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_92_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_93_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_94_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_95_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_96_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_97_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_98_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_99_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_100_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_101_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_102_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_103_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_104_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_105_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_106_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_107_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_108_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_109_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_110_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_111_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_112_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_113_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_114_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_115_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_116_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_117_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_118_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_119_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_120_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_121_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_122_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_123_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_124_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_125_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_126_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer2_out_127_blk_n);
    assign proc_5_data_PIPO_blk[0] = 1'b0;
    assign proc_5_start_FIFO_blk[0] = 1'b0 | (~myproject_U0.start_for_linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0_U.if_empty_n & myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.ap_idle & ~myproject_U0.start_for_linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0_U.if_write);
    assign proc_5_TLF_FIFO_blk[0] = 1'b0;
    assign proc_5_input_sync_blk[0] = 1'b0;
    assign proc_5_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_5[0] = dl_detect_out ? proc_dep_vld_vec_5_reg[0] : (proc_5_data_FIFO_blk[0] | proc_5_data_PIPO_blk[0] | proc_5_start_FIFO_blk[0] | proc_5_TLF_FIFO_blk[0] | proc_5_input_sync_blk[0] | proc_5_output_sync_blk[0]);
    assign proc_5_data_FIFO_blk[1] = 1'b0 | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_0_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_1_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_2_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_3_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_4_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_5_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_6_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_7_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_8_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_9_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_10_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_11_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_12_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_13_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_14_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_15_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_16_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_17_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_18_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_19_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_20_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_21_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_22_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_23_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_24_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_25_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_26_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_27_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_28_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_29_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_30_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_31_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_32_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_33_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_34_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_35_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_36_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_37_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_38_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_39_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_40_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_41_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_42_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_43_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_44_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_45_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_46_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_47_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_48_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_49_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_50_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_51_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_52_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_53_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_54_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_55_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_56_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_57_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_58_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_59_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_60_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_61_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_62_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_63_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_64_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_65_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_66_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_67_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_68_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_69_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_70_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_71_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_72_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_73_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_74_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_75_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_76_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_77_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_78_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_79_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_80_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_81_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_82_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_83_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_84_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_85_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_86_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_87_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_88_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_89_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_90_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_91_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_92_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_93_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_94_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_95_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_96_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_97_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_98_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_99_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_100_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_101_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_102_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_103_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_104_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_105_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_106_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_107_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_108_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_109_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_110_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_111_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_112_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_113_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_114_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_115_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_116_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_117_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_118_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_119_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_120_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_121_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_122_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_123_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_124_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_125_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_126_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.layer3_out_127_blk_n);
    assign proc_5_data_PIPO_blk[1] = 1'b0;
    assign proc_5_start_FIFO_blk[1] = 1'b0 | (~myproject_U0.start_for_clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0_U.if_full_n & myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.ap_start & ~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config3_U0.real_start & (trans_in_cnt_2 == trans_out_cnt_2) & ~myproject_U0.start_for_clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0_U.if_read);
    assign proc_5_TLF_FIFO_blk[1] = 1'b0;
    assign proc_5_input_sync_blk[1] = 1'b0;
    assign proc_5_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_5[1] = dl_detect_out ? proc_dep_vld_vec_5_reg[1] : (proc_5_data_FIFO_blk[1] | proc_5_data_PIPO_blk[1] | proc_5_start_FIFO_blk[1] | proc_5_TLF_FIFO_blk[1] | proc_5_input_sync_blk[1] | proc_5_output_sync_blk[1]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_5_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_5_reg <= proc_dep_vld_vec_5;
        end
    end
    assign in_chan_dep_vld_vec_5[0] = dep_chan_vld_4_5;
    assign in_chan_dep_data_vec_5[25 : 0] = dep_chan_data_4_5;
    assign token_in_vec_5[0] = token_4_5;
    assign in_chan_dep_vld_vec_5[1] = dep_chan_vld_6_5;
    assign in_chan_dep_data_vec_5[51 : 26] = dep_chan_data_6_5;
    assign token_in_vec_5[1] = token_6_5;
    assign dep_chan_vld_5_4 = out_chan_dep_vld_vec_5[0];
    assign dep_chan_data_5_4 = out_chan_dep_data_5;
    assign token_5_4 = token_out_vec_5[0];
    assign dep_chan_vld_5_6 = out_chan_dep_vld_vec_5[1];
    assign dep_chan_data_5_6 = out_chan_dep_data_5;
    assign token_5_6 = token_out_vec_5[1];

    // Process: myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0
    alveo_hls4ml_hls_deadlock_detect_unit #(26, 6, 3, 3) alveo_hls4ml_hls_deadlock_detect_unit_6 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_6),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_6),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_6),
        .token_in_vec(token_in_vec_6),
        .dl_detect_in(dl_detect_out),
        .origin(origin[6]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_6),
        .out_chan_dep_data(out_chan_dep_data_6),
        .token_out_vec(token_out_vec_6),
        .dl_detect_out(dl_in_vec[6]));

    assign proc_6_data_FIFO_blk[0] = 1'b0 | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_0_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_1_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_2_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_3_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_4_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_5_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_6_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_7_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_8_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_9_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_10_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_11_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_12_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_13_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_14_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_15_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_16_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_17_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_18_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_19_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_20_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_21_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_22_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_23_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_24_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_25_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_26_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_27_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_28_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_29_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_30_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_31_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_32_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_33_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_34_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_35_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_36_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_37_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_38_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_39_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_40_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_41_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_42_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_43_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_44_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_45_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_46_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_47_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_48_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_49_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_50_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_51_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_52_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_53_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_54_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_55_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_56_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_57_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_58_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_59_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_60_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_61_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_62_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_63_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_64_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_65_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_66_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_67_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_68_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_69_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_70_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_71_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_72_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_73_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_74_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_75_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_76_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_77_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_78_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_79_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_80_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_81_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_82_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_83_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_84_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_85_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_86_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_87_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_88_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_89_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_90_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_91_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_92_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_93_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_94_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_95_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_96_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_97_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_98_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_99_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_100_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_101_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_102_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_103_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_104_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_105_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_106_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_107_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_108_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_109_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_110_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_111_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_112_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_113_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_114_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_115_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_116_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_117_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_118_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_119_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_120_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_121_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_122_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_123_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_124_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_125_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_126_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer3_out_127_blk_n);
    assign proc_6_data_PIPO_blk[0] = 1'b0;
    assign proc_6_start_FIFO_blk[0] = 1'b0 | (~myproject_U0.start_for_clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0_U.if_empty_n & myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.ap_idle & ~myproject_U0.start_for_clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0_U.if_write);
    assign proc_6_TLF_FIFO_blk[0] = 1'b0;
    assign proc_6_input_sync_blk[0] = 1'b0;
    assign proc_6_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_6[0] = dl_detect_out ? proc_dep_vld_vec_6_reg[0] : (proc_6_data_FIFO_blk[0] | proc_6_data_PIPO_blk[0] | proc_6_start_FIFO_blk[0] | proc_6_TLF_FIFO_blk[0] | proc_6_input_sync_blk[0] | proc_6_output_sync_blk[0]);
    assign proc_6_data_FIFO_blk[1] = 1'b0 | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_0_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_1_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_2_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_3_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_4_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_5_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_6_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_7_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_8_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_9_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_10_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_11_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_12_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_13_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_14_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_15_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_16_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_17_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_18_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_19_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_20_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_21_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_22_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_23_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_24_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_25_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_26_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_27_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_28_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_29_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_30_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_31_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_32_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_33_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_34_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_35_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_36_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_37_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_38_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_39_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_40_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_41_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_42_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_43_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_44_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_45_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_46_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_47_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_48_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_49_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_50_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_51_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_52_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_53_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_54_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_55_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_56_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_57_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_58_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_59_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_60_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_61_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_62_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_63_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_64_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_65_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_66_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_67_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_68_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_69_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_70_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_71_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_72_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_73_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_74_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_75_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_76_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_77_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_78_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_79_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_80_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_81_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_82_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_83_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_84_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_85_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_86_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_87_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_88_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_89_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_90_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_91_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_92_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_93_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_94_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_95_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_96_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_97_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_98_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_99_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_100_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_101_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_102_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_103_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_104_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_105_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_106_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_107_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_108_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_109_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_110_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_111_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_112_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_113_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_114_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_115_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_116_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_117_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_118_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_119_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_120_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_121_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_122_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_123_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_124_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_125_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_126_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy1_127_blk_n);
    assign proc_6_data_PIPO_blk[1] = 1'b0;
    assign proc_6_start_FIFO_blk[1] = 1'b0 | (~myproject_U0.start_for_dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0_U.if_full_n & myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.ap_start & ~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.real_start & (trans_in_cnt_3 == trans_out_cnt_3) & ~myproject_U0.start_for_dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0_U.if_read);
    assign proc_6_TLF_FIFO_blk[1] = 1'b0;
    assign proc_6_input_sync_blk[1] = 1'b0;
    assign proc_6_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_6[1] = dl_detect_out ? proc_dep_vld_vec_6_reg[1] : (proc_6_data_FIFO_blk[1] | proc_6_data_PIPO_blk[1] | proc_6_start_FIFO_blk[1] | proc_6_TLF_FIFO_blk[1] | proc_6_input_sync_blk[1] | proc_6_output_sync_blk[1]);
    assign proc_6_data_FIFO_blk[2] = 1'b0 | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_0_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_1_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_2_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_3_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_4_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_5_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_6_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_7_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_8_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_9_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_10_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_11_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_12_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_13_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_14_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_15_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_16_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_17_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_18_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_19_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_20_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_21_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_22_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_23_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_24_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_25_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_26_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_27_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_28_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_29_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_30_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_31_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_32_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_33_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_34_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_35_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_36_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_37_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_38_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_39_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_40_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_41_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_42_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_43_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_44_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_45_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_46_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_47_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_48_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_49_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_50_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_51_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_52_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_53_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_54_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_55_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_56_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_57_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_58_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_59_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_60_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_61_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_62_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_63_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_64_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_65_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_66_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_67_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_68_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_69_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_70_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_71_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_72_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_73_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_74_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_75_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_76_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_77_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_78_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_79_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_80_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_81_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_82_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_83_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_84_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_85_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_86_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_87_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_88_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_89_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_90_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_91_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_92_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_93_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_94_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_95_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_96_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_97_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_98_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_99_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_100_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_101_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_102_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_103_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_104_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_105_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_106_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_107_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_108_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_109_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_110_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_111_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_112_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_113_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_114_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_115_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_116_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_117_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_118_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_119_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_120_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_121_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_122_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_123_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_124_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_125_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_126_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.layer28_cpy2_127_blk_n);
    assign proc_6_data_PIPO_blk[2] = 1'b0;
    assign proc_6_start_FIFO_blk[2] = 1'b0 | (~myproject_U0.start_for_dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0_U.if_full_n & myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.ap_start & ~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_128_U0.real_start & (trans_in_cnt_3 == trans_out_cnt_3) & ~myproject_U0.start_for_dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0_U.if_read);
    assign proc_6_TLF_FIFO_blk[2] = 1'b0;
    assign proc_6_input_sync_blk[2] = 1'b0;
    assign proc_6_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_6[2] = dl_detect_out ? proc_dep_vld_vec_6_reg[2] : (proc_6_data_FIFO_blk[2] | proc_6_data_PIPO_blk[2] | proc_6_start_FIFO_blk[2] | proc_6_TLF_FIFO_blk[2] | proc_6_input_sync_blk[2] | proc_6_output_sync_blk[2]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_6_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_6_reg <= proc_dep_vld_vec_6;
        end
    end
    assign in_chan_dep_vld_vec_6[0] = dep_chan_vld_5_6;
    assign in_chan_dep_data_vec_6[25 : 0] = dep_chan_data_5_6;
    assign token_in_vec_6[0] = token_5_6;
    assign in_chan_dep_vld_vec_6[1] = dep_chan_vld_7_6;
    assign in_chan_dep_data_vec_6[51 : 26] = dep_chan_data_7_6;
    assign token_in_vec_6[1] = token_7_6;
    assign in_chan_dep_vld_vec_6[2] = dep_chan_vld_8_6;
    assign in_chan_dep_data_vec_6[77 : 52] = dep_chan_data_8_6;
    assign token_in_vec_6[2] = token_8_6;
    assign dep_chan_vld_6_5 = out_chan_dep_vld_vec_6[0];
    assign dep_chan_data_6_5 = out_chan_dep_data_6;
    assign token_6_5 = token_out_vec_6[0];
    assign dep_chan_vld_6_7 = out_chan_dep_vld_vec_6[1];
    assign dep_chan_data_6_7 = out_chan_dep_data_6;
    assign token_6_7 = token_out_vec_6[1];
    assign dep_chan_vld_6_8 = out_chan_dep_vld_vec_6[2];
    assign dep_chan_data_6_8 = out_chan_dep_data_6;
    assign token_6_8 = token_out_vec_6[2];

    // Process: myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0
    alveo_hls4ml_hls_deadlock_detect_unit #(26, 7, 2, 2) alveo_hls4ml_hls_deadlock_detect_unit_7 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_7),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_7),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_7),
        .token_in_vec(token_in_vec_7),
        .dl_detect_in(dl_detect_out),
        .origin(origin[7]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_7),
        .out_chan_dep_data(out_chan_dep_data_7),
        .token_out_vec(token_out_vec_7),
        .dl_detect_out(dl_in_vec[7]));

    assign proc_7_data_FIFO_blk[0] = 1'b0 | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_0_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_1_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_2_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_3_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_4_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_5_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_6_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_7_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_8_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_9_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_10_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_11_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_12_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_13_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_14_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_15_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_16_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_17_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_18_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_19_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_20_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_21_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_22_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_23_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_24_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_25_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_26_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_27_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_28_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_29_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_30_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_31_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_32_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_33_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_34_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_35_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_36_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_37_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_38_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_39_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_40_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_41_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_42_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_43_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_44_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_45_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_46_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_47_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_48_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_49_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_50_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_51_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_52_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_53_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_54_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_55_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_56_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_57_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_58_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_59_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_60_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_61_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_62_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_63_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_64_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_65_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_66_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_67_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_68_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_69_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_70_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_71_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_72_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_73_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_74_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_75_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_76_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_77_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_78_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_79_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_80_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_81_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_82_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_83_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_84_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_85_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_86_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_87_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_88_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_89_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_90_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_91_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_92_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_93_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_94_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_95_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_96_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_97_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_98_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_99_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_100_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_101_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_102_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_103_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_104_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_105_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_106_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_107_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_108_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_109_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_110_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_111_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_112_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_113_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_114_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_115_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_116_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_117_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_118_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_119_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_120_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_121_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_122_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_123_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_124_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_125_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_126_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer28_cpy1_127_blk_n);
    assign proc_7_data_PIPO_blk[0] = 1'b0;
    assign proc_7_start_FIFO_blk[0] = 1'b0 | (~myproject_U0.start_for_dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0_U.if_empty_n & myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.ap_idle & ~myproject_U0.start_for_dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0_U.if_write);
    assign proc_7_TLF_FIFO_blk[0] = 1'b0;
    assign proc_7_input_sync_blk[0] = 1'b0;
    assign proc_7_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_7[0] = dl_detect_out ? proc_dep_vld_vec_7_reg[0] : (proc_7_data_FIFO_blk[0] | proc_7_data_PIPO_blk[0] | proc_7_start_FIFO_blk[0] | proc_7_TLF_FIFO_blk[0] | proc_7_input_sync_blk[0] | proc_7_output_sync_blk[0]);
    assign proc_7_data_FIFO_blk[1] = 1'b0 | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_0_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_1_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_2_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_3_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_4_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_5_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_6_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_7_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_8_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_9_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_10_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_11_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_12_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_13_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_14_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_15_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_16_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_17_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_18_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_19_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_20_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_21_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_22_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_23_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_24_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_25_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_26_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_27_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_28_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_29_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_30_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_31_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_32_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_33_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_34_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_35_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_36_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_37_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_38_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_39_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_40_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_41_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_42_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_43_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_44_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_45_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_46_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_47_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_48_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_49_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_50_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_51_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_52_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_53_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_54_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_55_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_56_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_57_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_58_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_59_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_60_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_61_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_62_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.layer4_out_63_blk_n);
    assign proc_7_data_PIPO_blk[1] = 1'b0;
    assign proc_7_start_FIFO_blk[1] = 1'b0 | (~myproject_U0.start_for_linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0_U.if_full_n & myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.ap_start & ~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config4_U0.real_start & (trans_in_cnt_4 == trans_out_cnt_4) & ~myproject_U0.start_for_linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0_U.if_read);
    assign proc_7_TLF_FIFO_blk[1] = 1'b0;
    assign proc_7_input_sync_blk[1] = 1'b0;
    assign proc_7_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_7[1] = dl_detect_out ? proc_dep_vld_vec_7_reg[1] : (proc_7_data_FIFO_blk[1] | proc_7_data_PIPO_blk[1] | proc_7_start_FIFO_blk[1] | proc_7_TLF_FIFO_blk[1] | proc_7_input_sync_blk[1] | proc_7_output_sync_blk[1]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_7_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_7_reg <= proc_dep_vld_vec_7;
        end
    end
    assign in_chan_dep_vld_vec_7[0] = dep_chan_vld_6_7;
    assign in_chan_dep_data_vec_7[25 : 0] = dep_chan_data_6_7;
    assign token_in_vec_7[0] = token_6_7;
    assign in_chan_dep_vld_vec_7[1] = dep_chan_vld_9_7;
    assign in_chan_dep_data_vec_7[51 : 26] = dep_chan_data_9_7;
    assign token_in_vec_7[1] = token_9_7;
    assign dep_chan_vld_7_6 = out_chan_dep_vld_vec_7[0];
    assign dep_chan_data_7_6 = out_chan_dep_data_7;
    assign token_7_6 = token_out_vec_7[0];
    assign dep_chan_vld_7_9 = out_chan_dep_vld_vec_7[1];
    assign dep_chan_data_7_9 = out_chan_dep_data_7;
    assign token_7_9 = token_out_vec_7[1];

    // Process: myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0
    alveo_hls4ml_hls_deadlock_detect_unit #(26, 8, 2, 2) alveo_hls4ml_hls_deadlock_detect_unit_8 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_8),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_8),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_8),
        .token_in_vec(token_in_vec_8),
        .dl_detect_in(dl_detect_out),
        .origin(origin[8]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_8),
        .out_chan_dep_data(out_chan_dep_data_8),
        .token_out_vec(token_out_vec_8),
        .dl_detect_out(dl_in_vec[8]));

    assign proc_8_data_FIFO_blk[0] = 1'b0 | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_0_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_1_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_2_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_3_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_4_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_5_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_6_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_7_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_8_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_9_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_10_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_11_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_12_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_13_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_14_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_15_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_16_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_17_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_18_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_19_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_20_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_21_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_22_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_23_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_24_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_25_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_26_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_27_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_28_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_29_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_30_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_31_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_32_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_33_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_34_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_35_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_36_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_37_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_38_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_39_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_40_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_41_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_42_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_43_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_44_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_45_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_46_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_47_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_48_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_49_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_50_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_51_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_52_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_53_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_54_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_55_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_56_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_57_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_58_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_59_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_60_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_61_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_62_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_63_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_64_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_65_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_66_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_67_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_68_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_69_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_70_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_71_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_72_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_73_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_74_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_75_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_76_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_77_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_78_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_79_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_80_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_81_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_82_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_83_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_84_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_85_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_86_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_87_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_88_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_89_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_90_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_91_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_92_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_93_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_94_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_95_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_96_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_97_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_98_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_99_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_100_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_101_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_102_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_103_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_104_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_105_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_106_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_107_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_108_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_109_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_110_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_111_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_112_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_113_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_114_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_115_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_116_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_117_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_118_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_119_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_120_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_121_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_122_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_123_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_124_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_125_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_126_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer28_cpy2_127_blk_n);
    assign proc_8_data_PIPO_blk[0] = 1'b0;
    assign proc_8_start_FIFO_blk[0] = 1'b0 | (~myproject_U0.start_for_dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0_U.if_empty_n & myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.ap_idle & ~myproject_U0.start_for_dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0_U.if_write);
    assign proc_8_TLF_FIFO_blk[0] = 1'b0;
    assign proc_8_input_sync_blk[0] = 1'b0;
    assign proc_8_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_8[0] = dl_detect_out ? proc_dep_vld_vec_8_reg[0] : (proc_8_data_FIFO_blk[0] | proc_8_data_PIPO_blk[0] | proc_8_start_FIFO_blk[0] | proc_8_TLF_FIFO_blk[0] | proc_8_input_sync_blk[0] | proc_8_output_sync_blk[0]);
    assign proc_8_data_FIFO_blk[1] = 1'b0 | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_0_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_1_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_2_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_3_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_4_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_5_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_6_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_7_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_8_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_9_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_10_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_11_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_12_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_13_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_14_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_15_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_16_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_17_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_18_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_19_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_20_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_21_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_22_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_23_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_24_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_25_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_26_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_27_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_28_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_29_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_30_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_31_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_32_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_33_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_34_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_35_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_36_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_37_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_38_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_39_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_40_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_41_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_42_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_43_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_44_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_45_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_46_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_47_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_48_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_49_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_50_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_51_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_52_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_53_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_54_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_55_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_56_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_57_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_58_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_59_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_60_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_61_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_62_blk_n) | (~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.layer6_out_63_blk_n);
    assign proc_8_data_PIPO_blk[1] = 1'b0;
    assign proc_8_start_FIFO_blk[1] = 1'b0 | (~myproject_U0.start_for_linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0_U.if_full_n & myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.ap_start & ~myproject_U0.dense_ap_fixed_16_6_5_3_0_ap_fixed_16_6_5_3_0_config6_U0.real_start & (trans_in_cnt_6 == trans_out_cnt_6) & ~myproject_U0.start_for_linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0_U.if_read);
    assign proc_8_TLF_FIFO_blk[1] = 1'b0;
    assign proc_8_input_sync_blk[1] = 1'b0;
    assign proc_8_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_8[1] = dl_detect_out ? proc_dep_vld_vec_8_reg[1] : (proc_8_data_FIFO_blk[1] | proc_8_data_PIPO_blk[1] | proc_8_start_FIFO_blk[1] | proc_8_TLF_FIFO_blk[1] | proc_8_input_sync_blk[1] | proc_8_output_sync_blk[1]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_8_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_8_reg <= proc_dep_vld_vec_8;
        end
    end
    assign in_chan_dep_vld_vec_8[0] = dep_chan_vld_6_8;
    assign in_chan_dep_data_vec_8[25 : 0] = dep_chan_data_6_8;
    assign token_in_vec_8[0] = token_6_8;
    assign in_chan_dep_vld_vec_8[1] = dep_chan_vld_11_8;
    assign in_chan_dep_data_vec_8[51 : 26] = dep_chan_data_11_8;
    assign token_in_vec_8[1] = token_11_8;
    assign dep_chan_vld_8_6 = out_chan_dep_vld_vec_8[0];
    assign dep_chan_data_8_6 = out_chan_dep_data_8;
    assign token_8_6 = token_out_vec_8[0];
    assign dep_chan_vld_8_11 = out_chan_dep_vld_vec_8[1];
    assign dep_chan_data_8_11 = out_chan_dep_data_8;
    assign token_8_11 = token_out_vec_8[1];

    // Process: myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0
    alveo_hls4ml_hls_deadlock_detect_unit #(26, 9, 2, 2) alveo_hls4ml_hls_deadlock_detect_unit_9 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_9),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_9),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_9),
        .token_in_vec(token_in_vec_9),
        .dl_detect_in(dl_detect_out),
        .origin(origin[9]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_9),
        .out_chan_dep_data(out_chan_dep_data_9),
        .token_out_vec(token_out_vec_9),
        .dl_detect_out(dl_in_vec[9]));

    assign proc_9_data_FIFO_blk[0] = 1'b0 | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_0_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_1_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_2_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_3_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_4_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_5_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_6_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_7_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_8_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_9_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_10_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_11_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_12_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_13_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_14_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_15_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_16_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_17_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_18_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_19_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_20_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_21_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_22_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_23_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_24_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_25_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_26_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_27_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_28_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_29_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_30_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_31_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_32_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_33_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_34_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_35_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_36_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_37_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_38_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_39_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_40_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_41_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_42_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_43_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_44_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_45_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_46_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_47_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_48_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_49_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_50_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_51_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_52_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_53_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_54_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_55_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_56_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_57_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_58_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_59_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_60_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_61_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_62_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer4_out_63_blk_n);
    assign proc_9_data_PIPO_blk[0] = 1'b0;
    assign proc_9_start_FIFO_blk[0] = 1'b0 | (~myproject_U0.start_for_linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0_U.if_empty_n & myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.ap_idle & ~myproject_U0.start_for_linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0_U.if_write);
    assign proc_9_TLF_FIFO_blk[0] = 1'b0;
    assign proc_9_input_sync_blk[0] = 1'b0;
    assign proc_9_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_9[0] = dl_detect_out ? proc_dep_vld_vec_9_reg[0] : (proc_9_data_FIFO_blk[0] | proc_9_data_PIPO_blk[0] | proc_9_start_FIFO_blk[0] | proc_9_TLF_FIFO_blk[0] | proc_9_input_sync_blk[0] | proc_9_output_sync_blk[0]);
    assign proc_9_data_FIFO_blk[1] = 1'b0 | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_0_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_1_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_2_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_3_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_4_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_5_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_6_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_7_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_8_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_9_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_10_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_11_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_12_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_13_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_14_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_15_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_16_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_17_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_18_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_19_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_20_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_21_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_22_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_23_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_24_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_25_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_26_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_27_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_28_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_29_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_30_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_31_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_32_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_33_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_34_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_35_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_36_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_37_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_38_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_39_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_40_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_41_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_42_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_43_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_44_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_45_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_46_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_47_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_48_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_49_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_50_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_51_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_52_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_53_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_54_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_55_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_56_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_57_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_58_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_59_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_60_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_61_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_62_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.layer8_out_63_blk_n);
    assign proc_9_data_PIPO_blk[1] = 1'b0;
    assign proc_9_start_FIFO_blk[1] = 1'b0 | (~myproject_U0.start_for_clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0_U.if_full_n & myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.ap_start & ~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config8_U0.real_start & (trans_in_cnt_5 == trans_out_cnt_5) & ~myproject_U0.start_for_clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0_U.if_read);
    assign proc_9_TLF_FIFO_blk[1] = 1'b0;
    assign proc_9_input_sync_blk[1] = 1'b0;
    assign proc_9_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_9[1] = dl_detect_out ? proc_dep_vld_vec_9_reg[1] : (proc_9_data_FIFO_blk[1] | proc_9_data_PIPO_blk[1] | proc_9_start_FIFO_blk[1] | proc_9_TLF_FIFO_blk[1] | proc_9_input_sync_blk[1] | proc_9_output_sync_blk[1]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_9_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_9_reg <= proc_dep_vld_vec_9;
        end
    end
    assign in_chan_dep_vld_vec_9[0] = dep_chan_vld_7_9;
    assign in_chan_dep_data_vec_9[25 : 0] = dep_chan_data_7_9;
    assign token_in_vec_9[0] = token_7_9;
    assign in_chan_dep_vld_vec_9[1] = dep_chan_vld_10_9;
    assign in_chan_dep_data_vec_9[51 : 26] = dep_chan_data_10_9;
    assign token_in_vec_9[1] = token_10_9;
    assign dep_chan_vld_9_7 = out_chan_dep_vld_vec_9[0];
    assign dep_chan_data_9_7 = out_chan_dep_data_9;
    assign token_9_7 = token_out_vec_9[0];
    assign dep_chan_vld_9_10 = out_chan_dep_vld_vec_9[1];
    assign dep_chan_data_9_10 = out_chan_dep_data_9;
    assign token_9_10 = token_out_vec_9[1];

    // Process: myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0
    alveo_hls4ml_hls_deadlock_detect_unit #(26, 10, 3, 3) alveo_hls4ml_hls_deadlock_detect_unit_10 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_10),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_10),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_10),
        .token_in_vec(token_in_vec_10),
        .dl_detect_in(dl_detect_out),
        .origin(origin[10]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_10),
        .out_chan_dep_data(out_chan_dep_data_10),
        .token_out_vec(token_out_vec_10),
        .dl_detect_out(dl_in_vec[10]));

    assign proc_10_data_FIFO_blk[0] = 1'b0 | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_0_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_1_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_2_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_3_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_4_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_5_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_6_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_7_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_8_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_9_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_10_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_11_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_12_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_13_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_14_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_15_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_16_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_17_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_18_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_19_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_20_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_21_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_22_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_23_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_24_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_25_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_26_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_27_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_28_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_29_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_30_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_31_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_32_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_33_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_34_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_35_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_36_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_37_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_38_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_39_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_40_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_41_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_42_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_43_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_44_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_45_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_46_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_47_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_48_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_49_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_50_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_51_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_52_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_53_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_54_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_55_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_56_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_57_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_58_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_59_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_60_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_61_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_62_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer8_out_63_blk_n);
    assign proc_10_data_PIPO_blk[0] = 1'b0;
    assign proc_10_start_FIFO_blk[0] = 1'b0 | (~myproject_U0.start_for_clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0_U.if_empty_n & myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.ap_idle & ~myproject_U0.start_for_clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0_U.if_write);
    assign proc_10_TLF_FIFO_blk[0] = 1'b0;
    assign proc_10_input_sync_blk[0] = 1'b0;
    assign proc_10_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_10[0] = dl_detect_out ? proc_dep_vld_vec_10_reg[0] : (proc_10_data_FIFO_blk[0] | proc_10_data_PIPO_blk[0] | proc_10_start_FIFO_blk[0] | proc_10_TLF_FIFO_blk[0] | proc_10_input_sync_blk[0] | proc_10_output_sync_blk[0]);
    assign proc_10_data_FIFO_blk[1] = 1'b0 | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_0_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_1_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_2_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_3_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_4_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_5_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_6_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_7_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_8_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_9_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_10_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_11_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_12_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_13_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_14_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_15_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_16_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_17_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_18_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_19_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_20_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_21_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_22_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_23_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_24_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_25_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_26_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_27_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_28_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_29_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_30_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_31_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_32_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_33_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_34_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_35_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_36_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_37_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_38_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_39_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_40_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_41_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_42_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_43_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_44_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_45_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_46_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_47_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_48_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_49_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_50_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_51_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_52_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_53_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_54_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_55_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_56_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_57_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_58_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_59_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_60_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_61_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_62_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy1_63_blk_n);
    assign proc_10_data_PIPO_blk[1] = 1'b0;
    assign proc_10_start_FIFO_blk[1] = 1'b0 | (~myproject_U0.start_for_srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0_U.if_full_n & myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.ap_start & ~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.real_start & (trans_in_cnt_8 == trans_out_cnt_8) & ~myproject_U0.start_for_srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0_U.if_read);
    assign proc_10_TLF_FIFO_blk[1] = 1'b0;
    assign proc_10_input_sync_blk[1] = 1'b0;
    assign proc_10_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_10[1] = dl_detect_out ? proc_dep_vld_vec_10_reg[1] : (proc_10_data_FIFO_blk[1] | proc_10_data_PIPO_blk[1] | proc_10_start_FIFO_blk[1] | proc_10_TLF_FIFO_blk[1] | proc_10_input_sync_blk[1] | proc_10_output_sync_blk[1]);
    assign proc_10_data_FIFO_blk[2] = 1'b0 | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_0_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_1_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_2_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_3_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_4_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_5_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_6_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_7_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_8_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_9_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_10_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_11_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_12_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_13_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_14_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_15_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_16_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_17_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_18_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_19_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_20_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_21_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_22_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_23_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_24_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_25_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_26_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_27_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_28_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_29_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_30_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_31_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_32_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_33_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_34_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_35_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_36_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_37_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_38_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_39_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_40_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_41_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_42_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_43_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_44_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_45_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_46_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_47_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_48_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_49_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_50_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_51_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_52_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_53_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_54_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_55_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_56_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_57_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_58_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_59_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_60_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_61_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_62_blk_n) | (~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.layer29_cpy2_63_blk_n);
    assign proc_10_data_PIPO_blk[2] = 1'b0;
    assign proc_10_start_FIFO_blk[2] = 1'b0 | (~myproject_U0.start_for_add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0_U.if_full_n & myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.ap_start & ~myproject_U0.clone_stream_ap_fixed_16_3_4_0_0_ap_fixed_32_16_5_3_0_64_U0.real_start & (trans_in_cnt_8 == trans_out_cnt_8) & ~myproject_U0.start_for_add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0_U.if_read);
    assign proc_10_TLF_FIFO_blk[2] = 1'b0;
    assign proc_10_input_sync_blk[2] = 1'b0;
    assign proc_10_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_10[2] = dl_detect_out ? proc_dep_vld_vec_10_reg[2] : (proc_10_data_FIFO_blk[2] | proc_10_data_PIPO_blk[2] | proc_10_start_FIFO_blk[2] | proc_10_TLF_FIFO_blk[2] | proc_10_input_sync_blk[2] | proc_10_output_sync_blk[2]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_10_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_10_reg <= proc_dep_vld_vec_10;
        end
    end
    assign in_chan_dep_vld_vec_10[0] = dep_chan_vld_9_10;
    assign in_chan_dep_data_vec_10[25 : 0] = dep_chan_data_9_10;
    assign token_in_vec_10[0] = token_9_10;
    assign in_chan_dep_vld_vec_10[1] = dep_chan_vld_13_10;
    assign in_chan_dep_data_vec_10[51 : 26] = dep_chan_data_13_10;
    assign token_in_vec_10[1] = token_13_10;
    assign in_chan_dep_vld_vec_10[2] = dep_chan_vld_18_10;
    assign in_chan_dep_data_vec_10[77 : 52] = dep_chan_data_18_10;
    assign token_in_vec_10[2] = token_18_10;
    assign dep_chan_vld_10_9 = out_chan_dep_vld_vec_10[0];
    assign dep_chan_data_10_9 = out_chan_dep_data_10;
    assign token_10_9 = token_out_vec_10[0];
    assign dep_chan_vld_10_13 = out_chan_dep_vld_vec_10[1];
    assign dep_chan_data_10_13 = out_chan_dep_data_10;
    assign token_10_13 = token_out_vec_10[1];
    assign dep_chan_vld_10_18 = out_chan_dep_vld_vec_10[2];
    assign dep_chan_data_10_18 = out_chan_dep_data_10;
    assign token_10_18 = token_out_vec_10[2];

    // Process: myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0
    alveo_hls4ml_hls_deadlock_detect_unit #(26, 11, 2, 2) alveo_hls4ml_hls_deadlock_detect_unit_11 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_11),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_11),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_11),
        .token_in_vec(token_in_vec_11),
        .dl_detect_in(dl_detect_out),
        .origin(origin[11]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_11),
        .out_chan_dep_data(out_chan_dep_data_11),
        .token_out_vec(token_out_vec_11),
        .dl_detect_out(dl_in_vec[11]));

    assign proc_11_data_FIFO_blk[0] = 1'b0 | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_0_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_1_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_2_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_3_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_4_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_5_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_6_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_7_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_8_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_9_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_10_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_11_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_12_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_13_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_14_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_15_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_16_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_17_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_18_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_19_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_20_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_21_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_22_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_23_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_24_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_25_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_26_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_27_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_28_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_29_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_30_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_31_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_32_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_33_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_34_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_35_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_36_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_37_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_38_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_39_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_40_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_41_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_42_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_43_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_44_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_45_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_46_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_47_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_48_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_49_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_50_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_51_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_52_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_53_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_54_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_55_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_56_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_57_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_58_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_59_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_60_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_61_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_62_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer6_out_63_blk_n);
    assign proc_11_data_PIPO_blk[0] = 1'b0;
    assign proc_11_start_FIFO_blk[0] = 1'b0 | (~myproject_U0.start_for_linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0_U.if_empty_n & myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.ap_idle & ~myproject_U0.start_for_linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0_U.if_write);
    assign proc_11_TLF_FIFO_blk[0] = 1'b0;
    assign proc_11_input_sync_blk[0] = 1'b0;
    assign proc_11_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_11[0] = dl_detect_out ? proc_dep_vld_vec_11_reg[0] : (proc_11_data_FIFO_blk[0] | proc_11_data_PIPO_blk[0] | proc_11_start_FIFO_blk[0] | proc_11_TLF_FIFO_blk[0] | proc_11_input_sync_blk[0] | proc_11_output_sync_blk[0]);
    assign proc_11_data_FIFO_blk[1] = 1'b0 | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_0_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_1_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_2_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_3_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_4_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_5_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_6_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_7_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_8_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_9_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_10_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_11_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_12_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_13_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_14_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_15_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_16_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_17_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_18_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_19_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_20_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_21_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_22_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_23_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_24_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_25_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_26_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_27_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_28_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_29_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_30_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_31_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_32_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_33_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_34_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_35_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_36_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_37_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_38_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_39_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_40_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_41_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_42_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_43_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_44_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_45_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_46_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_47_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_48_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_49_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_50_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_51_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_52_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_53_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_54_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_55_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_56_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_57_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_58_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_59_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_60_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_61_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_62_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.layer9_out_63_blk_n);
    assign proc_11_data_PIPO_blk[1] = 1'b0;
    assign proc_11_start_FIFO_blk[1] = 1'b0 | (~myproject_U0.start_for_explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0_U.if_full_n & myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.ap_start & ~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_10_3_4_0_0_linear_config9_U0.real_start & (trans_in_cnt_7 == trans_out_cnt_7) & ~myproject_U0.start_for_explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0_U.if_read);
    assign proc_11_TLF_FIFO_blk[1] = 1'b0;
    assign proc_11_input_sync_blk[1] = 1'b0;
    assign proc_11_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_11[1] = dl_detect_out ? proc_dep_vld_vec_11_reg[1] : (proc_11_data_FIFO_blk[1] | proc_11_data_PIPO_blk[1] | proc_11_start_FIFO_blk[1] | proc_11_TLF_FIFO_blk[1] | proc_11_input_sync_blk[1] | proc_11_output_sync_blk[1]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_11_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_11_reg <= proc_dep_vld_vec_11;
        end
    end
    assign in_chan_dep_vld_vec_11[0] = dep_chan_vld_8_11;
    assign in_chan_dep_data_vec_11[25 : 0] = dep_chan_data_8_11;
    assign token_in_vec_11[0] = token_8_11;
    assign in_chan_dep_vld_vec_11[1] = dep_chan_vld_12_11;
    assign in_chan_dep_data_vec_11[51 : 26] = dep_chan_data_12_11;
    assign token_in_vec_11[1] = token_12_11;
    assign dep_chan_vld_11_8 = out_chan_dep_vld_vec_11[0];
    assign dep_chan_data_11_8 = out_chan_dep_data_11;
    assign token_11_8 = token_out_vec_11[0];
    assign dep_chan_vld_11_12 = out_chan_dep_vld_vec_11[1];
    assign dep_chan_data_11_12 = out_chan_dep_data_11;
    assign token_11_12 = token_out_vec_11[1];

    // Process: myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0
    alveo_hls4ml_hls_deadlock_detect_unit #(26, 12, 2, 2) alveo_hls4ml_hls_deadlock_detect_unit_12 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_12),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_12),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_12),
        .token_in_vec(token_in_vec_12),
        .dl_detect_in(dl_detect_out),
        .origin(origin[12]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_12),
        .out_chan_dep_data(out_chan_dep_data_12),
        .token_out_vec(token_out_vec_12),
        .dl_detect_out(dl_in_vec[12]));

    assign proc_12_data_FIFO_blk[0] = 1'b0 | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_0_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_1_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_2_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_3_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_4_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_5_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_6_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_7_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_8_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_9_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_10_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_11_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_12_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_13_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_14_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_15_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_16_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_17_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_18_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_19_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_20_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_21_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_22_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_23_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_24_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_25_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_26_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_27_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_28_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_29_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_30_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_31_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_32_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_33_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_34_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_35_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_36_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_37_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_38_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_39_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_40_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_41_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_42_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_43_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_44_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_45_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_46_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_47_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_48_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_49_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_50_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_51_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_52_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_53_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_54_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_55_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_56_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_57_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_58_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_59_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_60_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_61_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_62_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer9_out_63_blk_n);
    assign proc_12_data_PIPO_blk[0] = 1'b0;
    assign proc_12_start_FIFO_blk[0] = 1'b0 | (~myproject_U0.start_for_explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0_U.if_empty_n & myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.ap_idle & ~myproject_U0.start_for_explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0_U.if_write);
    assign proc_12_TLF_FIFO_blk[0] = 1'b0;
    assign proc_12_input_sync_blk[0] = 1'b0;
    assign proc_12_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_12[0] = dl_detect_out ? proc_dep_vld_vec_12_reg[0] : (proc_12_data_FIFO_blk[0] | proc_12_data_PIPO_blk[0] | proc_12_start_FIFO_blk[0] | proc_12_TLF_FIFO_blk[0] | proc_12_input_sync_blk[0] | proc_12_output_sync_blk[0]);
    assign proc_12_data_FIFO_blk[1] = 1'b0 | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_0_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_1_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_2_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_3_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_4_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_5_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_6_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_7_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_8_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_9_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_10_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_11_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_12_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_13_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_14_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_15_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_16_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_17_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_18_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_19_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_20_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_21_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_22_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_23_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_24_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_25_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_26_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_27_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_28_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_29_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_30_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_31_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_32_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_33_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_34_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_35_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_36_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_37_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_38_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_39_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_40_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_41_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_42_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_43_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_44_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_45_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_46_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_47_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_48_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_49_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_50_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_51_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_52_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_53_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_54_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_55_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_56_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_57_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_58_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_59_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_60_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_61_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_62_blk_n) | (~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.layer10_out_63_blk_n);
    assign proc_12_data_PIPO_blk[1] = 1'b0;
    assign proc_12_start_FIFO_blk[1] = 1'b0 | (~myproject_U0.start_for_linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0_U.if_full_n & myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.ap_start & ~myproject_U0.explogvar_ap_fixed_10_3_4_0_0_ap_fixed_16_6_5_3_0_config10_U0.real_start & (trans_in_cnt_9 == trans_out_cnt_9) & ~myproject_U0.start_for_linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0_U.if_read);
    assign proc_12_TLF_FIFO_blk[1] = 1'b0;
    assign proc_12_input_sync_blk[1] = 1'b0;
    assign proc_12_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_12[1] = dl_detect_out ? proc_dep_vld_vec_12_reg[1] : (proc_12_data_FIFO_blk[1] | proc_12_data_PIPO_blk[1] | proc_12_start_FIFO_blk[1] | proc_12_TLF_FIFO_blk[1] | proc_12_input_sync_blk[1] | proc_12_output_sync_blk[1]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_12_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_12_reg <= proc_dep_vld_vec_12;
        end
    end
    assign in_chan_dep_vld_vec_12[0] = dep_chan_vld_11_12;
    assign in_chan_dep_data_vec_12[25 : 0] = dep_chan_data_11_12;
    assign token_in_vec_12[0] = token_11_12;
    assign in_chan_dep_vld_vec_12[1] = dep_chan_vld_14_12;
    assign in_chan_dep_data_vec_12[51 : 26] = dep_chan_data_14_12;
    assign token_in_vec_12[1] = token_14_12;
    assign dep_chan_vld_12_11 = out_chan_dep_vld_vec_12[0];
    assign dep_chan_data_12_11 = out_chan_dep_data_12;
    assign token_12_11 = token_out_vec_12[0];
    assign dep_chan_vld_12_14 = out_chan_dep_vld_vec_12[1];
    assign dep_chan_data_12_14 = out_chan_dep_data_12;
    assign token_12_14 = token_out_vec_12[1];

    // Process: myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0
    alveo_hls4ml_hls_deadlock_detect_unit #(26, 13, 2, 2) alveo_hls4ml_hls_deadlock_detect_unit_13 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_13),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_13),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_13),
        .token_in_vec(token_in_vec_13),
        .dl_detect_in(dl_detect_out),
        .origin(origin[13]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_13),
        .out_chan_dep_data(out_chan_dep_data_13),
        .token_out_vec(token_out_vec_13),
        .dl_detect_out(dl_in_vec[13]));

    assign proc_13_data_FIFO_blk[0] = 1'b0 | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_0_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_1_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_2_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_3_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_4_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_5_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_6_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_7_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_8_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_9_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_10_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_11_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_12_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_13_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_14_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_15_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_16_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_17_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_18_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_19_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_20_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_21_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_22_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_23_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_24_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_25_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_26_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_27_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_28_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_29_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_30_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_31_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_32_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_33_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_34_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_35_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_36_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_37_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_38_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_39_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_40_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_41_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_42_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_43_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_44_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_45_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_46_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_47_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_48_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_49_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_50_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_51_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_52_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_53_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_54_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_55_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_56_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_57_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_58_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_59_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_60_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_61_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_62_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer29_cpy1_63_blk_n);
    assign proc_13_data_PIPO_blk[0] = 1'b0;
    assign proc_13_start_FIFO_blk[0] = 1'b0 | (~myproject_U0.start_for_srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0_U.if_empty_n & myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.ap_idle & ~myproject_U0.start_for_srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0_U.if_write);
    assign proc_13_TLF_FIFO_blk[0] = 1'b0;
    assign proc_13_input_sync_blk[0] = 1'b0;
    assign proc_13_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_13[0] = dl_detect_out ? proc_dep_vld_vec_13_reg[0] : (proc_13_data_FIFO_blk[0] | proc_13_data_PIPO_blk[0] | proc_13_start_FIFO_blk[0] | proc_13_TLF_FIFO_blk[0] | proc_13_input_sync_blk[0] | proc_13_output_sync_blk[0]);
    assign proc_13_data_FIFO_blk[1] = 1'b0 | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_0_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_1_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_2_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_3_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_4_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_5_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_6_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_7_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_8_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_9_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_10_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_11_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_12_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_13_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_14_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_15_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_16_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_17_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_18_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_19_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_20_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_21_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_22_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_23_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_24_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_25_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_26_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_27_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_28_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_29_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_30_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_31_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_32_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_33_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_34_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_35_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_36_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_37_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_38_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_39_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_40_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_41_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_42_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_43_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_44_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_45_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_46_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_47_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_48_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_49_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_50_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_51_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_52_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_53_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_54_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_55_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_56_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_57_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_58_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_59_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_60_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_61_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_62_blk_n) | (~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.layer11_out_63_blk_n);
    assign proc_13_data_PIPO_blk[1] = 1'b0;
    assign proc_13_start_FIFO_blk[1] = 1'b0 | (~myproject_U0.start_for_linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0_U.if_full_n & myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.ap_start & ~myproject_U0.srn_ap_fixed_32_16_5_3_0_ap_fixed_32_16_5_3_0_config11_U0.real_start & (trans_in_cnt_10 == trans_out_cnt_10) & ~myproject_U0.start_for_linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0_U.if_read);
    assign proc_13_TLF_FIFO_blk[1] = 1'b0;
    assign proc_13_input_sync_blk[1] = 1'b0;
    assign proc_13_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_13[1] = dl_detect_out ? proc_dep_vld_vec_13_reg[1] : (proc_13_data_FIFO_blk[1] | proc_13_data_PIPO_blk[1] | proc_13_start_FIFO_blk[1] | proc_13_TLF_FIFO_blk[1] | proc_13_input_sync_blk[1] | proc_13_output_sync_blk[1]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_13_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_13_reg <= proc_dep_vld_vec_13;
        end
    end
    assign in_chan_dep_vld_vec_13[0] = dep_chan_vld_10_13;
    assign in_chan_dep_data_vec_13[25 : 0] = dep_chan_data_10_13;
    assign token_in_vec_13[0] = token_10_13;
    assign in_chan_dep_vld_vec_13[1] = dep_chan_vld_15_13;
    assign in_chan_dep_data_vec_13[51 : 26] = dep_chan_data_15_13;
    assign token_in_vec_13[1] = token_15_13;
    assign dep_chan_vld_13_10 = out_chan_dep_vld_vec_13[0];
    assign dep_chan_data_13_10 = out_chan_dep_data_13;
    assign token_13_10 = token_out_vec_13[0];
    assign dep_chan_vld_13_15 = out_chan_dep_vld_vec_13[1];
    assign dep_chan_data_13_15 = out_chan_dep_data_13;
    assign token_13_15 = token_out_vec_13[1];

    // Process: myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0
    alveo_hls4ml_hls_deadlock_detect_unit #(26, 14, 2, 2) alveo_hls4ml_hls_deadlock_detect_unit_14 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_14),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_14),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_14),
        .token_in_vec(token_in_vec_14),
        .dl_detect_in(dl_detect_out),
        .origin(origin[14]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_14),
        .out_chan_dep_data(out_chan_dep_data_14),
        .token_out_vec(token_out_vec_14),
        .dl_detect_out(dl_in_vec[14]));

    assign proc_14_data_FIFO_blk[0] = 1'b0 | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_0_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_1_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_2_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_3_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_4_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_5_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_6_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_7_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_8_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_9_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_10_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_11_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_12_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_13_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_14_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_15_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_16_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_17_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_18_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_19_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_20_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_21_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_22_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_23_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_24_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_25_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_26_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_27_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_28_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_29_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_30_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_31_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_32_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_33_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_34_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_35_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_36_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_37_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_38_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_39_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_40_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_41_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_42_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_43_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_44_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_45_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_46_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_47_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_48_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_49_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_50_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_51_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_52_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_53_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_54_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_55_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_56_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_57_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_58_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_59_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_60_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_61_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_62_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer10_out_63_blk_n);
    assign proc_14_data_PIPO_blk[0] = 1'b0;
    assign proc_14_start_FIFO_blk[0] = 1'b0 | (~myproject_U0.start_for_linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0_U.if_empty_n & myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.ap_idle & ~myproject_U0.start_for_linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0_U.if_write);
    assign proc_14_TLF_FIFO_blk[0] = 1'b0;
    assign proc_14_input_sync_blk[0] = 1'b0;
    assign proc_14_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_14[0] = dl_detect_out ? proc_dep_vld_vec_14_reg[0] : (proc_14_data_FIFO_blk[0] | proc_14_data_PIPO_blk[0] | proc_14_start_FIFO_blk[0] | proc_14_TLF_FIFO_blk[0] | proc_14_input_sync_blk[0] | proc_14_output_sync_blk[0]);
    assign proc_14_data_FIFO_blk[1] = 1'b0 | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_0_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_1_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_2_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_3_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_4_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_5_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_6_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_7_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_8_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_9_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_10_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_11_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_12_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_13_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_14_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_15_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_16_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_17_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_18_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_19_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_20_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_21_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_22_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_23_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_24_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_25_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_26_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_27_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_28_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_29_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_30_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_31_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_32_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_33_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_34_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_35_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_36_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_37_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_38_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_39_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_40_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_41_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_42_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_43_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_44_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_45_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_46_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_47_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_48_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_49_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_50_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_51_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_52_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_53_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_54_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_55_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_56_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_57_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_58_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_59_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_60_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_61_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_62_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.layer12_out_63_blk_n);
    assign proc_14_data_PIPO_blk[1] = 1'b0;
    assign proc_14_start_FIFO_blk[1] = 1'b0 | (~myproject_U0.start_for_multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0_U.if_full_n & myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.ap_start & ~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_18_8_4_0_0_linear_config12_U0.real_start & (trans_in_cnt_11 == trans_out_cnt_11) & ~myproject_U0.start_for_multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0_U.if_read);
    assign proc_14_TLF_FIFO_blk[1] = 1'b0;
    assign proc_14_input_sync_blk[1] = 1'b0;
    assign proc_14_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_14[1] = dl_detect_out ? proc_dep_vld_vec_14_reg[1] : (proc_14_data_FIFO_blk[1] | proc_14_data_PIPO_blk[1] | proc_14_start_FIFO_blk[1] | proc_14_TLF_FIFO_blk[1] | proc_14_input_sync_blk[1] | proc_14_output_sync_blk[1]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_14_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_14_reg <= proc_dep_vld_vec_14;
        end
    end
    assign in_chan_dep_vld_vec_14[0] = dep_chan_vld_12_14;
    assign in_chan_dep_data_vec_14[25 : 0] = dep_chan_data_12_14;
    assign token_in_vec_14[0] = token_12_14;
    assign in_chan_dep_vld_vec_14[1] = dep_chan_vld_16_14;
    assign in_chan_dep_data_vec_14[51 : 26] = dep_chan_data_16_14;
    assign token_in_vec_14[1] = token_16_14;
    assign dep_chan_vld_14_12 = out_chan_dep_vld_vec_14[0];
    assign dep_chan_data_14_12 = out_chan_dep_data_14;
    assign token_14_12 = token_out_vec_14[0];
    assign dep_chan_vld_14_16 = out_chan_dep_vld_vec_14[1];
    assign dep_chan_data_14_16 = out_chan_dep_data_14;
    assign token_14_16 = token_out_vec_14[1];

    // Process: myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0
    alveo_hls4ml_hls_deadlock_detect_unit #(26, 15, 2, 2) alveo_hls4ml_hls_deadlock_detect_unit_15 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_15),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_15),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_15),
        .token_in_vec(token_in_vec_15),
        .dl_detect_in(dl_detect_out),
        .origin(origin[15]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_15),
        .out_chan_dep_data(out_chan_dep_data_15),
        .token_out_vec(token_out_vec_15),
        .dl_detect_out(dl_in_vec[15]));

    assign proc_15_data_FIFO_blk[0] = 1'b0 | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_0_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_1_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_2_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_3_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_4_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_5_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_6_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_7_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_8_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_9_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_10_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_11_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_12_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_13_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_14_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_15_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_16_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_17_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_18_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_19_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_20_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_21_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_22_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_23_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_24_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_25_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_26_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_27_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_28_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_29_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_30_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_31_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_32_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_33_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_34_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_35_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_36_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_37_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_38_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_39_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_40_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_41_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_42_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_43_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_44_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_45_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_46_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_47_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_48_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_49_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_50_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_51_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_52_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_53_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_54_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_55_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_56_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_57_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_58_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_59_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_60_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_61_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_62_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer11_out_63_blk_n);
    assign proc_15_data_PIPO_blk[0] = 1'b0;
    assign proc_15_start_FIFO_blk[0] = 1'b0 | (~myproject_U0.start_for_linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0_U.if_empty_n & myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.ap_idle & ~myproject_U0.start_for_linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0_U.if_write);
    assign proc_15_TLF_FIFO_blk[0] = 1'b0;
    assign proc_15_input_sync_blk[0] = 1'b0;
    assign proc_15_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_15[0] = dl_detect_out ? proc_dep_vld_vec_15_reg[0] : (proc_15_data_FIFO_blk[0] | proc_15_data_PIPO_blk[0] | proc_15_start_FIFO_blk[0] | proc_15_TLF_FIFO_blk[0] | proc_15_input_sync_blk[0] | proc_15_output_sync_blk[0]);
    assign proc_15_data_FIFO_blk[1] = 1'b0 | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_0_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_1_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_2_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_3_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_4_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_5_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_6_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_7_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_8_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_9_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_10_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_11_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_12_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_13_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_14_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_15_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_16_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_17_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_18_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_19_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_20_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_21_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_22_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_23_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_24_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_25_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_26_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_27_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_28_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_29_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_30_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_31_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_32_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_33_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_34_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_35_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_36_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_37_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_38_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_39_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_40_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_41_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_42_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_43_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_44_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_45_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_46_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_47_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_48_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_49_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_50_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_51_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_52_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_53_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_54_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_55_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_56_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_57_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_58_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_59_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_60_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_61_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_62_blk_n) | (~myproject_U0.linear_ap_fixed_32_16_5_3_0_ap_fixed_16_3_4_0_0_linear_config13_U0.layer13_out_63_blk_n);
    assign proc_15_data_PIPO_blk[1] = 1'b0;
    assign proc_15_start_FIFO_blk[1] = 1'b0;
    assign proc_15_TLF_FIFO_blk[1] = 1'b0;
    assign proc_15_input_sync_blk[1] = 1'b0;
    assign proc_15_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_15[1] = dl_detect_out ? proc_dep_vld_vec_15_reg[1] : (proc_15_data_FIFO_blk[1] | proc_15_data_PIPO_blk[1] | proc_15_start_FIFO_blk[1] | proc_15_TLF_FIFO_blk[1] | proc_15_input_sync_blk[1] | proc_15_output_sync_blk[1]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_15_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_15_reg <= proc_dep_vld_vec_15;
        end
    end
    assign in_chan_dep_vld_vec_15[0] = dep_chan_vld_13_15;
    assign in_chan_dep_data_vec_15[25 : 0] = dep_chan_data_13_15;
    assign token_in_vec_15[0] = token_13_15;
    assign in_chan_dep_vld_vec_15[1] = dep_chan_vld_16_15;
    assign in_chan_dep_data_vec_15[51 : 26] = dep_chan_data_16_15;
    assign token_in_vec_15[1] = token_16_15;
    assign dep_chan_vld_15_13 = out_chan_dep_vld_vec_15[0];
    assign dep_chan_data_15_13 = out_chan_dep_data_15;
    assign token_15_13 = token_out_vec_15[0];
    assign dep_chan_vld_15_16 = out_chan_dep_vld_vec_15[1];
    assign dep_chan_data_15_16 = out_chan_dep_data_15;
    assign token_15_16 = token_out_vec_15[1];

    // Process: myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0
    alveo_hls4ml_hls_deadlock_detect_unit #(26, 16, 3, 3) alveo_hls4ml_hls_deadlock_detect_unit_16 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_16),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_16),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_16),
        .token_in_vec(token_in_vec_16),
        .dl_detect_in(dl_detect_out),
        .origin(origin[16]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_16),
        .out_chan_dep_data(out_chan_dep_data_16),
        .token_out_vec(token_out_vec_16),
        .dl_detect_out(dl_in_vec[16]));

    assign proc_16_data_FIFO_blk[0] = 1'b0 | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_0_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_1_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_2_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_3_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_4_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_5_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_6_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_7_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_8_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_9_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_10_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_11_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_12_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_13_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_14_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_15_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_16_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_17_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_18_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_19_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_20_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_21_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_22_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_23_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_24_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_25_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_26_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_27_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_28_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_29_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_30_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_31_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_32_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_33_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_34_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_35_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_36_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_37_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_38_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_39_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_40_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_41_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_42_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_43_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_44_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_45_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_46_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_47_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_48_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_49_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_50_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_51_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_52_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_53_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_54_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_55_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_56_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_57_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_58_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_59_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_60_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_61_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_62_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer12_out_63_blk_n);
    assign proc_16_data_PIPO_blk[0] = 1'b0;
    assign proc_16_start_FIFO_blk[0] = 1'b0 | (~myproject_U0.start_for_multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0_U.if_empty_n & myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.ap_idle & ~myproject_U0.start_for_multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0_U.if_write);
    assign proc_16_TLF_FIFO_blk[0] = 1'b0;
    assign proc_16_input_sync_blk[0] = 1'b0;
    assign proc_16_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_16[0] = dl_detect_out ? proc_dep_vld_vec_16_reg[0] : (proc_16_data_FIFO_blk[0] | proc_16_data_PIPO_blk[0] | proc_16_start_FIFO_blk[0] | proc_16_TLF_FIFO_blk[0] | proc_16_input_sync_blk[0] | proc_16_output_sync_blk[0]);
    assign proc_16_data_FIFO_blk[1] = 1'b0 | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_0_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_1_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_2_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_3_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_4_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_5_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_6_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_7_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_8_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_9_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_10_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_11_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_12_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_13_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_14_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_15_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_16_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_17_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_18_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_19_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_20_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_21_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_22_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_23_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_24_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_25_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_26_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_27_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_28_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_29_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_30_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_31_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_32_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_33_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_34_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_35_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_36_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_37_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_38_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_39_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_40_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_41_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_42_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_43_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_44_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_45_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_46_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_47_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_48_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_49_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_50_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_51_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_52_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_53_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_54_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_55_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_56_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_57_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_58_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_59_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_60_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_61_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_62_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer13_out_63_blk_n);
    assign proc_16_data_PIPO_blk[1] = 1'b0;
    assign proc_16_start_FIFO_blk[1] = 1'b0;
    assign proc_16_TLF_FIFO_blk[1] = 1'b0;
    assign proc_16_input_sync_blk[1] = 1'b0;
    assign proc_16_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_16[1] = dl_detect_out ? proc_dep_vld_vec_16_reg[1] : (proc_16_data_FIFO_blk[1] | proc_16_data_PIPO_blk[1] | proc_16_start_FIFO_blk[1] | proc_16_TLF_FIFO_blk[1] | proc_16_input_sync_blk[1] | proc_16_output_sync_blk[1]);
    assign proc_16_data_FIFO_blk[2] = 1'b0 | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_0_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_1_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_2_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_3_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_4_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_5_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_6_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_7_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_8_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_9_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_10_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_11_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_12_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_13_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_14_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_15_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_16_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_17_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_18_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_19_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_20_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_21_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_22_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_23_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_24_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_25_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_26_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_27_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_28_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_29_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_30_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_31_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_32_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_33_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_34_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_35_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_36_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_37_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_38_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_39_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_40_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_41_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_42_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_43_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_44_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_45_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_46_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_47_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_48_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_49_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_50_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_51_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_52_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_53_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_54_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_55_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_56_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_57_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_58_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_59_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_60_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_61_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_62_blk_n) | (~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.layer14_out_63_blk_n);
    assign proc_16_data_PIPO_blk[2] = 1'b0;
    assign proc_16_start_FIFO_blk[2] = 1'b0 | (~myproject_U0.start_for_linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0_U.if_full_n & myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.ap_start & ~myproject_U0.multiply_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config14_U0.real_start & (trans_in_cnt_12 == trans_out_cnt_12) & ~myproject_U0.start_for_linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0_U.if_read);
    assign proc_16_TLF_FIFO_blk[2] = 1'b0;
    assign proc_16_input_sync_blk[2] = 1'b0;
    assign proc_16_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_16[2] = dl_detect_out ? proc_dep_vld_vec_16_reg[2] : (proc_16_data_FIFO_blk[2] | proc_16_data_PIPO_blk[2] | proc_16_start_FIFO_blk[2] | proc_16_TLF_FIFO_blk[2] | proc_16_input_sync_blk[2] | proc_16_output_sync_blk[2]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_16_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_16_reg <= proc_dep_vld_vec_16;
        end
    end
    assign in_chan_dep_vld_vec_16[0] = dep_chan_vld_14_16;
    assign in_chan_dep_data_vec_16[25 : 0] = dep_chan_data_14_16;
    assign token_in_vec_16[0] = token_14_16;
    assign in_chan_dep_vld_vec_16[1] = dep_chan_vld_15_16;
    assign in_chan_dep_data_vec_16[51 : 26] = dep_chan_data_15_16;
    assign token_in_vec_16[1] = token_15_16;
    assign in_chan_dep_vld_vec_16[2] = dep_chan_vld_17_16;
    assign in_chan_dep_data_vec_16[77 : 52] = dep_chan_data_17_16;
    assign token_in_vec_16[2] = token_17_16;
    assign dep_chan_vld_16_14 = out_chan_dep_vld_vec_16[0];
    assign dep_chan_data_16_14 = out_chan_dep_data_16;
    assign token_16_14 = token_out_vec_16[0];
    assign dep_chan_vld_16_15 = out_chan_dep_vld_vec_16[1];
    assign dep_chan_data_16_15 = out_chan_dep_data_16;
    assign token_16_15 = token_out_vec_16[1];
    assign dep_chan_vld_16_17 = out_chan_dep_vld_vec_16[2];
    assign dep_chan_data_16_17 = out_chan_dep_data_16;
    assign token_16_17 = token_out_vec_16[2];

    // Process: myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0
    alveo_hls4ml_hls_deadlock_detect_unit #(26, 17, 2, 2) alveo_hls4ml_hls_deadlock_detect_unit_17 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_17),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_17),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_17),
        .token_in_vec(token_in_vec_17),
        .dl_detect_in(dl_detect_out),
        .origin(origin[17]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_17),
        .out_chan_dep_data(out_chan_dep_data_17),
        .token_out_vec(token_out_vec_17),
        .dl_detect_out(dl_in_vec[17]));

    assign proc_17_data_FIFO_blk[0] = 1'b0 | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_0_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_1_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_2_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_3_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_4_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_5_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_6_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_7_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_8_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_9_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_10_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_11_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_12_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_13_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_14_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_15_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_16_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_17_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_18_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_19_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_20_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_21_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_22_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_23_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_24_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_25_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_26_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_27_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_28_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_29_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_30_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_31_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_32_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_33_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_34_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_35_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_36_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_37_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_38_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_39_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_40_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_41_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_42_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_43_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_44_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_45_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_46_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_47_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_48_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_49_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_50_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_51_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_52_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_53_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_54_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_55_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_56_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_57_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_58_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_59_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_60_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_61_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_62_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer14_out_63_blk_n);
    assign proc_17_data_PIPO_blk[0] = 1'b0;
    assign proc_17_start_FIFO_blk[0] = 1'b0 | (~myproject_U0.start_for_linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0_U.if_empty_n & myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.ap_idle & ~myproject_U0.start_for_linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0_U.if_write);
    assign proc_17_TLF_FIFO_blk[0] = 1'b0;
    assign proc_17_input_sync_blk[0] = 1'b0;
    assign proc_17_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_17[0] = dl_detect_out ? proc_dep_vld_vec_17_reg[0] : (proc_17_data_FIFO_blk[0] | proc_17_data_PIPO_blk[0] | proc_17_start_FIFO_blk[0] | proc_17_TLF_FIFO_blk[0] | proc_17_input_sync_blk[0] | proc_17_output_sync_blk[0]);
    assign proc_17_data_FIFO_blk[1] = 1'b0 | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_0_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_1_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_2_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_3_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_4_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_5_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_6_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_7_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_8_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_9_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_10_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_11_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_12_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_13_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_14_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_15_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_16_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_17_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_18_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_19_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_20_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_21_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_22_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_23_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_24_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_25_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_26_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_27_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_28_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_29_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_30_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_31_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_32_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_33_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_34_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_35_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_36_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_37_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_38_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_39_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_40_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_41_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_42_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_43_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_44_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_45_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_46_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_47_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_48_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_49_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_50_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_51_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_52_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_53_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_54_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_55_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_56_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_57_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_58_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_59_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_60_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_61_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_62_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config15_U0.layer15_out_63_blk_n);
    assign proc_17_data_PIPO_blk[1] = 1'b0;
    assign proc_17_start_FIFO_blk[1] = 1'b0;
    assign proc_17_TLF_FIFO_blk[1] = 1'b0;
    assign proc_17_input_sync_blk[1] = 1'b0;
    assign proc_17_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_17[1] = dl_detect_out ? proc_dep_vld_vec_17_reg[1] : (proc_17_data_FIFO_blk[1] | proc_17_data_PIPO_blk[1] | proc_17_start_FIFO_blk[1] | proc_17_TLF_FIFO_blk[1] | proc_17_input_sync_blk[1] | proc_17_output_sync_blk[1]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_17_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_17_reg <= proc_dep_vld_vec_17;
        end
    end
    assign in_chan_dep_vld_vec_17[0] = dep_chan_vld_16_17;
    assign in_chan_dep_data_vec_17[25 : 0] = dep_chan_data_16_17;
    assign token_in_vec_17[0] = token_16_17;
    assign in_chan_dep_vld_vec_17[1] = dep_chan_vld_18_17;
    assign in_chan_dep_data_vec_17[51 : 26] = dep_chan_data_18_17;
    assign token_in_vec_17[1] = token_18_17;
    assign dep_chan_vld_17_16 = out_chan_dep_vld_vec_17[0];
    assign dep_chan_data_17_16 = out_chan_dep_data_17;
    assign token_17_16 = token_out_vec_17[0];
    assign dep_chan_vld_17_18 = out_chan_dep_vld_vec_17[1];
    assign dep_chan_data_17_18 = out_chan_dep_data_17;
    assign token_17_18 = token_out_vec_17[1];

    // Process: myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0
    alveo_hls4ml_hls_deadlock_detect_unit #(26, 18, 3, 3) alveo_hls4ml_hls_deadlock_detect_unit_18 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_18),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_18),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_18),
        .token_in_vec(token_in_vec_18),
        .dl_detect_in(dl_detect_out),
        .origin(origin[18]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_18),
        .out_chan_dep_data(out_chan_dep_data_18),
        .token_out_vec(token_out_vec_18),
        .dl_detect_out(dl_in_vec[18]));

    assign proc_18_data_FIFO_blk[0] = 1'b0 | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_0_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_1_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_2_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_3_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_4_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_5_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_6_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_7_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_8_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_9_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_10_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_11_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_12_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_13_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_14_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_15_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_16_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_17_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_18_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_19_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_20_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_21_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_22_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_23_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_24_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_25_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_26_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_27_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_28_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_29_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_30_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_31_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_32_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_33_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_34_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_35_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_36_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_37_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_38_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_39_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_40_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_41_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_42_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_43_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_44_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_45_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_46_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_47_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_48_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_49_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_50_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_51_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_52_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_53_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_54_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_55_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_56_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_57_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_58_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_59_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_60_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_61_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_62_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer29_cpy2_63_blk_n);
    assign proc_18_data_PIPO_blk[0] = 1'b0;
    assign proc_18_start_FIFO_blk[0] = 1'b0 | (~myproject_U0.start_for_add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0_U.if_empty_n & myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.ap_idle & ~myproject_U0.start_for_add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0_U.if_write);
    assign proc_18_TLF_FIFO_blk[0] = 1'b0;
    assign proc_18_input_sync_blk[0] = 1'b0;
    assign proc_18_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_18[0] = dl_detect_out ? proc_dep_vld_vec_18_reg[0] : (proc_18_data_FIFO_blk[0] | proc_18_data_PIPO_blk[0] | proc_18_start_FIFO_blk[0] | proc_18_TLF_FIFO_blk[0] | proc_18_input_sync_blk[0] | proc_18_output_sync_blk[0]);
    assign proc_18_data_FIFO_blk[1] = 1'b0 | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_0_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_1_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_2_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_3_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_4_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_5_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_6_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_7_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_8_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_9_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_10_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_11_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_12_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_13_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_14_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_15_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_16_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_17_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_18_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_19_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_20_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_21_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_22_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_23_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_24_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_25_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_26_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_27_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_28_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_29_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_30_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_31_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_32_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_33_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_34_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_35_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_36_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_37_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_38_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_39_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_40_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_41_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_42_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_43_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_44_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_45_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_46_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_47_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_48_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_49_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_50_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_51_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_52_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_53_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_54_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_55_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_56_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_57_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_58_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_59_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_60_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_61_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_62_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer15_out_63_blk_n);
    assign proc_18_data_PIPO_blk[1] = 1'b0;
    assign proc_18_start_FIFO_blk[1] = 1'b0;
    assign proc_18_TLF_FIFO_blk[1] = 1'b0;
    assign proc_18_input_sync_blk[1] = 1'b0;
    assign proc_18_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_18[1] = dl_detect_out ? proc_dep_vld_vec_18_reg[1] : (proc_18_data_FIFO_blk[1] | proc_18_data_PIPO_blk[1] | proc_18_start_FIFO_blk[1] | proc_18_TLF_FIFO_blk[1] | proc_18_input_sync_blk[1] | proc_18_output_sync_blk[1]);
    assign proc_18_data_FIFO_blk[2] = 1'b0 | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_0_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_1_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_2_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_3_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_4_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_5_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_6_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_7_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_8_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_9_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_10_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_11_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_12_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_13_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_14_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_15_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_16_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_17_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_18_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_19_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_20_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_21_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_22_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_23_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_24_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_25_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_26_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_27_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_28_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_29_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_30_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_31_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_32_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_33_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_34_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_35_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_36_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_37_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_38_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_39_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_40_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_41_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_42_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_43_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_44_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_45_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_46_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_47_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_48_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_49_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_50_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_51_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_52_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_53_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_54_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_55_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_56_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_57_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_58_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_59_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_60_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_61_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_62_blk_n) | (~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.layer16_out_63_blk_n);
    assign proc_18_data_PIPO_blk[2] = 1'b0;
    assign proc_18_start_FIFO_blk[2] = 1'b0 | (~myproject_U0.start_for_linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0_U.if_full_n & myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.ap_start & ~myproject_U0.add_ap_fixed_ap_fixed_16_3_4_0_0_ap_fixed_16_6_5_3_0_config16_U0.real_start & (trans_in_cnt_13 == trans_out_cnt_13) & ~myproject_U0.start_for_linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0_U.if_read);
    assign proc_18_TLF_FIFO_blk[2] = 1'b0;
    assign proc_18_input_sync_blk[2] = 1'b0;
    assign proc_18_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_18[2] = dl_detect_out ? proc_dep_vld_vec_18_reg[2] : (proc_18_data_FIFO_blk[2] | proc_18_data_PIPO_blk[2] | proc_18_start_FIFO_blk[2] | proc_18_TLF_FIFO_blk[2] | proc_18_input_sync_blk[2] | proc_18_output_sync_blk[2]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_18_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_18_reg <= proc_dep_vld_vec_18;
        end
    end
    assign in_chan_dep_vld_vec_18[0] = dep_chan_vld_10_18;
    assign in_chan_dep_data_vec_18[25 : 0] = dep_chan_data_10_18;
    assign token_in_vec_18[0] = token_10_18;
    assign in_chan_dep_vld_vec_18[1] = dep_chan_vld_17_18;
    assign in_chan_dep_data_vec_18[51 : 26] = dep_chan_data_17_18;
    assign token_in_vec_18[1] = token_17_18;
    assign in_chan_dep_vld_vec_18[2] = dep_chan_vld_19_18;
    assign in_chan_dep_data_vec_18[77 : 52] = dep_chan_data_19_18;
    assign token_in_vec_18[2] = token_19_18;
    assign dep_chan_vld_18_10 = out_chan_dep_vld_vec_18[0];
    assign dep_chan_data_18_10 = out_chan_dep_data_18;
    assign token_18_10 = token_out_vec_18[0];
    assign dep_chan_vld_18_17 = out_chan_dep_vld_vec_18[1];
    assign dep_chan_data_18_17 = out_chan_dep_data_18;
    assign token_18_17 = token_out_vec_18[1];
    assign dep_chan_vld_18_19 = out_chan_dep_vld_vec_18[2];
    assign dep_chan_data_18_19 = out_chan_dep_data_18;
    assign token_18_19 = token_out_vec_18[2];

    // Process: myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0
    alveo_hls4ml_hls_deadlock_detect_unit #(26, 19, 2, 2) alveo_hls4ml_hls_deadlock_detect_unit_19 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_19),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_19),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_19),
        .token_in_vec(token_in_vec_19),
        .dl_detect_in(dl_detect_out),
        .origin(origin[19]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_19),
        .out_chan_dep_data(out_chan_dep_data_19),
        .token_out_vec(token_out_vec_19),
        .dl_detect_out(dl_in_vec[19]));

    assign proc_19_data_FIFO_blk[0] = 1'b0 | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_0_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_1_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_2_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_3_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_4_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_5_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_6_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_7_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_8_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_9_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_10_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_11_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_12_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_13_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_14_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_15_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_16_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_17_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_18_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_19_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_20_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_21_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_22_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_23_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_24_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_25_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_26_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_27_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_28_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_29_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_30_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_31_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_32_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_33_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_34_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_35_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_36_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_37_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_38_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_39_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_40_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_41_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_42_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_43_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_44_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_45_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_46_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_47_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_48_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_49_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_50_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_51_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_52_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_53_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_54_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_55_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_56_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_57_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_58_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_59_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_60_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_61_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_62_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer16_out_63_blk_n);
    assign proc_19_data_PIPO_blk[0] = 1'b0;
    assign proc_19_start_FIFO_blk[0] = 1'b0 | (~myproject_U0.start_for_linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0_U.if_empty_n & myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.ap_idle & ~myproject_U0.start_for_linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0_U.if_write);
    assign proc_19_TLF_FIFO_blk[0] = 1'b0;
    assign proc_19_input_sync_blk[0] = 1'b0;
    assign proc_19_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_19[0] = dl_detect_out ? proc_dep_vld_vec_19_reg[0] : (proc_19_data_FIFO_blk[0] | proc_19_data_PIPO_blk[0] | proc_19_start_FIFO_blk[0] | proc_19_TLF_FIFO_blk[0] | proc_19_input_sync_blk[0] | proc_19_output_sync_blk[0]);
    assign proc_19_data_FIFO_blk[1] = 1'b0 | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_0_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_1_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_2_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_3_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_4_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_5_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_6_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_7_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_8_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_9_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_10_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_11_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_12_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_13_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_14_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_15_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_16_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_17_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_18_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_19_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_20_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_21_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_22_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_23_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_24_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_25_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_26_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_27_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_28_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_29_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_30_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_31_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_32_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_33_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_34_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_35_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_36_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_37_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_38_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_39_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_40_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_41_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_42_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_43_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_44_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_45_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_46_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_47_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_48_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_49_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_50_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_51_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_52_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_53_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_54_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_55_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_56_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_57_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_58_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_59_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_60_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_61_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_62_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.layer18_out_63_blk_n);
    assign proc_19_data_PIPO_blk[1] = 1'b0;
    assign proc_19_start_FIFO_blk[1] = 1'b0 | (~myproject_U0.start_for_gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0_U.if_full_n & myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.ap_start & ~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config18_U0.real_start & (trans_in_cnt_14 == trans_out_cnt_14) & ~myproject_U0.start_for_gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0_U.if_read);
    assign proc_19_TLF_FIFO_blk[1] = 1'b0;
    assign proc_19_input_sync_blk[1] = 1'b0;
    assign proc_19_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_19[1] = dl_detect_out ? proc_dep_vld_vec_19_reg[1] : (proc_19_data_FIFO_blk[1] | proc_19_data_PIPO_blk[1] | proc_19_start_FIFO_blk[1] | proc_19_TLF_FIFO_blk[1] | proc_19_input_sync_blk[1] | proc_19_output_sync_blk[1]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_19_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_19_reg <= proc_dep_vld_vec_19;
        end
    end
    assign in_chan_dep_vld_vec_19[0] = dep_chan_vld_18_19;
    assign in_chan_dep_data_vec_19[25 : 0] = dep_chan_data_18_19;
    assign token_in_vec_19[0] = token_18_19;
    assign in_chan_dep_vld_vec_19[1] = dep_chan_vld_20_19;
    assign in_chan_dep_data_vec_19[51 : 26] = dep_chan_data_20_19;
    assign token_in_vec_19[1] = token_20_19;
    assign dep_chan_vld_19_18 = out_chan_dep_vld_vec_19[0];
    assign dep_chan_data_19_18 = out_chan_dep_data_19;
    assign token_19_18 = token_out_vec_19[0];
    assign dep_chan_vld_19_20 = out_chan_dep_vld_vec_19[1];
    assign dep_chan_data_19_20 = out_chan_dep_data_19;
    assign token_19_20 = token_out_vec_19[1];

    // Process: myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0
    alveo_hls4ml_hls_deadlock_detect_unit #(26, 20, 3, 3) alveo_hls4ml_hls_deadlock_detect_unit_20 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_20),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_20),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_20),
        .token_in_vec(token_in_vec_20),
        .dl_detect_in(dl_detect_out),
        .origin(origin[20]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_20),
        .out_chan_dep_data(out_chan_dep_data_20),
        .token_out_vec(token_out_vec_20),
        .dl_detect_out(dl_in_vec[20]));

    assign proc_20_data_FIFO_blk[0] = 1'b0 | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_0_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_1_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_2_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_3_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_4_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_5_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_6_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_7_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_8_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_9_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_10_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_11_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_12_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_13_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_14_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_15_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_16_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_17_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_18_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_19_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_20_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_21_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_22_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_23_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_24_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_25_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_26_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_27_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_28_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_29_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_30_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_31_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_32_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_33_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_34_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_35_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_36_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_37_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_38_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_39_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_40_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_41_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_42_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_43_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_44_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_45_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_46_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_47_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_48_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_49_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_50_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_51_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_52_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_53_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_54_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_55_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_56_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_57_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_58_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_59_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_60_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_61_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_62_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.in_stream2_63_blk_n);
    assign proc_20_data_PIPO_blk[0] = 1'b0;
    assign proc_20_start_FIFO_blk[0] = 1'b0;
    assign proc_20_TLF_FIFO_blk[0] = 1'b0;
    assign proc_20_input_sync_blk[0] = 1'b0;
    assign proc_20_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_20[0] = dl_detect_out ? proc_dep_vld_vec_20_reg[0] : (proc_20_data_FIFO_blk[0] | proc_20_data_PIPO_blk[0] | proc_20_start_FIFO_blk[0] | proc_20_TLF_FIFO_blk[0] | proc_20_input_sync_blk[0] | proc_20_output_sync_blk[0]);
    assign proc_20_data_FIFO_blk[1] = 1'b0 | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_0_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_1_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_2_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_3_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_4_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_5_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_6_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_7_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_8_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_9_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_10_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_11_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_12_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_13_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_14_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_15_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_16_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_17_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_18_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_19_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_20_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_21_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_22_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_23_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_24_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_25_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_26_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_27_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_28_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_29_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_30_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_31_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_32_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_33_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_34_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_35_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_36_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_37_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_38_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_39_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_40_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_41_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_42_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_43_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_44_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_45_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_46_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_47_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_48_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_49_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_50_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_51_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_52_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_53_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_54_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_55_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_56_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_57_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_58_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_59_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_60_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_61_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_62_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer18_out_63_blk_n);
    assign proc_20_data_PIPO_blk[1] = 1'b0;
    assign proc_20_start_FIFO_blk[1] = 1'b0 | (~myproject_U0.start_for_gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0_U.if_empty_n & myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.ap_idle & ~myproject_U0.start_for_gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0_U.if_write);
    assign proc_20_TLF_FIFO_blk[1] = 1'b0;
    assign proc_20_input_sync_blk[1] = 1'b0;
    assign proc_20_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_20[1] = dl_detect_out ? proc_dep_vld_vec_20_reg[1] : (proc_20_data_FIFO_blk[1] | proc_20_data_PIPO_blk[1] | proc_20_start_FIFO_blk[1] | proc_20_TLF_FIFO_blk[1] | proc_20_input_sync_blk[1] | proc_20_output_sync_blk[1]);
    assign proc_20_data_FIFO_blk[2] = 1'b0 | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_0_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_1_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_2_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_3_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_4_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_5_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_6_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_7_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_8_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_9_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_10_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_11_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_12_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_13_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_14_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_15_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_16_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_17_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_18_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_19_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_20_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_21_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_22_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_23_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_24_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_25_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_26_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_27_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_28_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_29_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_30_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_31_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_32_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_33_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_34_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_35_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_36_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_37_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_38_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_39_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_40_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_41_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_42_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_43_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_44_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_45_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_46_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_47_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_48_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_49_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_50_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_51_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_52_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_53_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_54_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_55_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_56_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_57_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_58_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_59_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_60_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_61_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_62_blk_n) | (~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.layer19_out_63_blk_n);
    assign proc_20_data_PIPO_blk[2] = 1'b0;
    assign proc_20_start_FIFO_blk[2] = 1'b0 | (~myproject_U0.start_for_linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0_U.if_full_n & myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.ap_start & ~myproject_U0.gru_stack_array_ap_fixed_ap_fixed_ap_fixed_33_4_5_3_0_config19_U0.real_start & (trans_in_cnt_15 == trans_out_cnt_15) & ~myproject_U0.start_for_linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0_U.if_read);
    assign proc_20_TLF_FIFO_blk[2] = 1'b0;
    assign proc_20_input_sync_blk[2] = 1'b0;
    assign proc_20_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_20[2] = dl_detect_out ? proc_dep_vld_vec_20_reg[2] : (proc_20_data_FIFO_blk[2] | proc_20_data_PIPO_blk[2] | proc_20_start_FIFO_blk[2] | proc_20_TLF_FIFO_blk[2] | proc_20_input_sync_blk[2] | proc_20_output_sync_blk[2]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_20_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_20_reg <= proc_dep_vld_vec_20;
        end
    end
    assign in_chan_dep_vld_vec_20[0] = dep_chan_vld_2_20;
    assign in_chan_dep_data_vec_20[25 : 0] = dep_chan_data_2_20;
    assign token_in_vec_20[0] = token_2_20;
    assign in_chan_dep_vld_vec_20[1] = dep_chan_vld_19_20;
    assign in_chan_dep_data_vec_20[51 : 26] = dep_chan_data_19_20;
    assign token_in_vec_20[1] = token_19_20;
    assign in_chan_dep_vld_vec_20[2] = dep_chan_vld_21_20;
    assign in_chan_dep_data_vec_20[77 : 52] = dep_chan_data_21_20;
    assign token_in_vec_20[2] = token_21_20;
    assign dep_chan_vld_20_2 = out_chan_dep_vld_vec_20[0];
    assign dep_chan_data_20_2 = out_chan_dep_data_20;
    assign token_20_2 = token_out_vec_20[0];
    assign dep_chan_vld_20_19 = out_chan_dep_vld_vec_20[1];
    assign dep_chan_data_20_19 = out_chan_dep_data_20;
    assign token_20_19 = token_out_vec_20[1];
    assign dep_chan_vld_20_21 = out_chan_dep_vld_vec_20[2];
    assign dep_chan_data_20_21 = out_chan_dep_data_20;
    assign token_20_21 = token_out_vec_20[2];

    // Process: myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0
    alveo_hls4ml_hls_deadlock_detect_unit #(26, 21, 2, 2) alveo_hls4ml_hls_deadlock_detect_unit_21 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_21),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_21),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_21),
        .token_in_vec(token_in_vec_21),
        .dl_detect_in(dl_detect_out),
        .origin(origin[21]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_21),
        .out_chan_dep_data(out_chan_dep_data_21),
        .token_out_vec(token_out_vec_21),
        .dl_detect_out(dl_in_vec[21]));

    assign proc_21_data_FIFO_blk[0] = 1'b0 | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_0_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_1_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_2_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_3_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_4_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_5_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_6_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_7_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_8_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_9_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_10_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_11_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_12_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_13_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_14_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_15_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_16_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_17_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_18_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_19_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_20_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_21_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_22_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_23_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_24_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_25_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_26_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_27_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_28_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_29_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_30_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_31_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_32_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_33_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_34_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_35_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_36_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_37_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_38_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_39_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_40_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_41_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_42_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_43_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_44_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_45_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_46_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_47_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_48_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_49_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_50_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_51_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_52_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_53_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_54_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_55_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_56_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_57_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_58_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_59_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_60_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_61_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_62_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer19_out_63_blk_n);
    assign proc_21_data_PIPO_blk[0] = 1'b0;
    assign proc_21_start_FIFO_blk[0] = 1'b0 | (~myproject_U0.start_for_linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0_U.if_empty_n & myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.ap_idle & ~myproject_U0.start_for_linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0_U.if_write);
    assign proc_21_TLF_FIFO_blk[0] = 1'b0;
    assign proc_21_input_sync_blk[0] = 1'b0;
    assign proc_21_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_21[0] = dl_detect_out ? proc_dep_vld_vec_21_reg[0] : (proc_21_data_FIFO_blk[0] | proc_21_data_PIPO_blk[0] | proc_21_start_FIFO_blk[0] | proc_21_TLF_FIFO_blk[0] | proc_21_input_sync_blk[0] | proc_21_output_sync_blk[0]);
    assign proc_21_data_FIFO_blk[1] = 1'b0 | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_0_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_1_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_2_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_3_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_4_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_5_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_6_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_7_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_8_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_9_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_10_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_11_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_12_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_13_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_14_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_15_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_16_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_17_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_18_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_19_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_20_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_21_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_22_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_23_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_24_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_25_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_26_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_27_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_28_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_29_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_30_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_31_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_32_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_33_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_34_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_35_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_36_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_37_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_38_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_39_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_40_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_41_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_42_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_43_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_44_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_45_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_46_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_47_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_48_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_49_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_50_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_51_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_52_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_53_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_54_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_55_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_56_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_57_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_58_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_59_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_60_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_61_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_62_blk_n) | (~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.layer20_out_63_blk_n);
    assign proc_21_data_PIPO_blk[1] = 1'b0;
    assign proc_21_start_FIFO_blk[1] = 1'b0 | (~myproject_U0.start_for_pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0_U.if_full_n & myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.ap_start & ~myproject_U0.linear_ap_fixed_33_4_5_3_0_ap_fixed_16_3_4_0_0_linear_config20_U0.real_start & (trans_in_cnt_16 == trans_out_cnt_16) & ~myproject_U0.start_for_pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0_U.if_read);
    assign proc_21_TLF_FIFO_blk[1] = 1'b0;
    assign proc_21_input_sync_blk[1] = 1'b0;
    assign proc_21_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_21[1] = dl_detect_out ? proc_dep_vld_vec_21_reg[1] : (proc_21_data_FIFO_blk[1] | proc_21_data_PIPO_blk[1] | proc_21_start_FIFO_blk[1] | proc_21_TLF_FIFO_blk[1] | proc_21_input_sync_blk[1] | proc_21_output_sync_blk[1]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_21_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_21_reg <= proc_dep_vld_vec_21;
        end
    end
    assign in_chan_dep_vld_vec_21[0] = dep_chan_vld_20_21;
    assign in_chan_dep_data_vec_21[25 : 0] = dep_chan_data_20_21;
    assign token_in_vec_21[0] = token_20_21;
    assign in_chan_dep_vld_vec_21[1] = dep_chan_vld_22_21;
    assign in_chan_dep_data_vec_21[51 : 26] = dep_chan_data_22_21;
    assign token_in_vec_21[1] = token_22_21;
    assign dep_chan_vld_21_20 = out_chan_dep_vld_vec_21[0];
    assign dep_chan_data_21_20 = out_chan_dep_data_21;
    assign token_21_20 = token_out_vec_21[0];
    assign dep_chan_vld_21_22 = out_chan_dep_vld_vec_21[1];
    assign dep_chan_data_21_22 = out_chan_dep_data_21;
    assign token_21_22 = token_out_vec_21[1];

    // Process: myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0
    alveo_hls4ml_hls_deadlock_detect_unit #(26, 22, 2, 2) alveo_hls4ml_hls_deadlock_detect_unit_22 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_22),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_22),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_22),
        .token_in_vec(token_in_vec_22),
        .dl_detect_in(dl_detect_out),
        .origin(origin[22]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_22),
        .out_chan_dep_data(out_chan_dep_data_22),
        .token_out_vec(token_out_vec_22),
        .dl_detect_out(dl_in_vec[22]));

    assign proc_22_data_FIFO_blk[0] = 1'b0 | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_0_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_1_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_2_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_3_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_4_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_5_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_6_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_7_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_8_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_9_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_10_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_11_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_12_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_13_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_14_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_15_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_16_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_17_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_18_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_19_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_20_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_21_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_22_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_23_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_24_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_25_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_26_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_27_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_28_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_29_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_30_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_31_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_32_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_33_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_34_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_35_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_36_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_37_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_38_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_39_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_40_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_41_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_42_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_43_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_44_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_45_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_46_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_47_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_48_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_49_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_50_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_51_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_52_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_53_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_54_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_55_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_56_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_57_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_58_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_59_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_60_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_61_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_62_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer20_out_63_blk_n);
    assign proc_22_data_PIPO_blk[0] = 1'b0;
    assign proc_22_start_FIFO_blk[0] = 1'b0 | (~myproject_U0.start_for_pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0_U.if_empty_n & myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.ap_idle & ~myproject_U0.start_for_pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0_U.if_write);
    assign proc_22_TLF_FIFO_blk[0] = 1'b0;
    assign proc_22_input_sync_blk[0] = 1'b0;
    assign proc_22_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_22[0] = dl_detect_out ? proc_dep_vld_vec_22_reg[0] : (proc_22_data_FIFO_blk[0] | proc_22_data_PIPO_blk[0] | proc_22_start_FIFO_blk[0] | proc_22_TLF_FIFO_blk[0] | proc_22_input_sync_blk[0] | proc_22_output_sync_blk[0]);
    assign proc_22_data_FIFO_blk[1] = 1'b0 | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer26_out_0_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer26_out_1_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer26_out_2_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.layer26_out_3_blk_n);
    assign proc_22_data_PIPO_blk[1] = 1'b0;
    assign proc_22_start_FIFO_blk[1] = 1'b0 | (~myproject_U0.start_for_linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config23_U0_U.if_full_n & myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.ap_start & ~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config26_U0.real_start & (trans_in_cnt_17 == trans_out_cnt_17) & ~myproject_U0.start_for_linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config23_U0_U.if_read);
    assign proc_22_TLF_FIFO_blk[1] = 1'b0;
    assign proc_22_input_sync_blk[1] = 1'b0;
    assign proc_22_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_22[1] = dl_detect_out ? proc_dep_vld_vec_22_reg[1] : (proc_22_data_FIFO_blk[1] | proc_22_data_PIPO_blk[1] | proc_22_start_FIFO_blk[1] | proc_22_TLF_FIFO_blk[1] | proc_22_input_sync_blk[1] | proc_22_output_sync_blk[1]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_22_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_22_reg <= proc_dep_vld_vec_22;
        end
    end
    assign in_chan_dep_vld_vec_22[0] = dep_chan_vld_21_22;
    assign in_chan_dep_data_vec_22[25 : 0] = dep_chan_data_21_22;
    assign token_in_vec_22[0] = token_21_22;
    assign in_chan_dep_vld_vec_22[1] = dep_chan_vld_23_22;
    assign in_chan_dep_data_vec_22[51 : 26] = dep_chan_data_23_22;
    assign token_in_vec_22[1] = token_23_22;
    assign dep_chan_vld_22_21 = out_chan_dep_vld_vec_22[0];
    assign dep_chan_data_22_21 = out_chan_dep_data_22;
    assign token_22_21 = token_out_vec_22[0];
    assign dep_chan_vld_22_23 = out_chan_dep_vld_vec_22[1];
    assign dep_chan_data_22_23 = out_chan_dep_data_22;
    assign token_22_23 = token_out_vec_22[1];

    // Process: myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config23_U0
    alveo_hls4ml_hls_deadlock_detect_unit #(26, 23, 2, 2) alveo_hls4ml_hls_deadlock_detect_unit_23 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_23),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_23),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_23),
        .token_in_vec(token_in_vec_23),
        .dl_detect_in(dl_detect_out),
        .origin(origin[23]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_23),
        .out_chan_dep_data(out_chan_dep_data_23),
        .token_out_vec(token_out_vec_23),
        .dl_detect_out(dl_in_vec[23]));

    assign proc_23_data_FIFO_blk[0] = 1'b0 | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config23_U0.layer26_out_0_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config23_U0.layer26_out_1_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config23_U0.layer26_out_2_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config23_U0.layer26_out_3_blk_n);
    assign proc_23_data_PIPO_blk[0] = 1'b0;
    assign proc_23_start_FIFO_blk[0] = 1'b0 | (~myproject_U0.start_for_linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config23_U0_U.if_empty_n & myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config23_U0.ap_idle & ~myproject_U0.start_for_linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config23_U0_U.if_write);
    assign proc_23_TLF_FIFO_blk[0] = 1'b0;
    assign proc_23_input_sync_blk[0] = 1'b0;
    assign proc_23_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_23[0] = dl_detect_out ? proc_dep_vld_vec_23_reg[0] : (proc_23_data_FIFO_blk[0] | proc_23_data_PIPO_blk[0] | proc_23_start_FIFO_blk[0] | proc_23_TLF_FIFO_blk[0] | proc_23_input_sync_blk[0] | proc_23_output_sync_blk[0]);
    assign proc_23_data_FIFO_blk[1] = 1'b0 | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config23_U0.layer23_out_0_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config23_U0.layer23_out_1_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config23_U0.layer23_out_2_blk_n) | (~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config23_U0.layer23_out_3_blk_n);
    assign proc_23_data_PIPO_blk[1] = 1'b0;
    assign proc_23_start_FIFO_blk[1] = 1'b0 | (~myproject_U0.start_for_pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0_U.if_full_n & myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config23_U0.ap_start & ~myproject_U0.linear_ap_fixed_16_6_5_3_0_ap_fixed_16_3_4_0_0_linear_config23_U0.real_start & (trans_in_cnt_18 == trans_out_cnt_18) & ~myproject_U0.start_for_pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0_U.if_read);
    assign proc_23_TLF_FIFO_blk[1] = 1'b0;
    assign proc_23_input_sync_blk[1] = 1'b0;
    assign proc_23_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_23[1] = dl_detect_out ? proc_dep_vld_vec_23_reg[1] : (proc_23_data_FIFO_blk[1] | proc_23_data_PIPO_blk[1] | proc_23_start_FIFO_blk[1] | proc_23_TLF_FIFO_blk[1] | proc_23_input_sync_blk[1] | proc_23_output_sync_blk[1]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_23_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_23_reg <= proc_dep_vld_vec_23;
        end
    end
    assign in_chan_dep_vld_vec_23[0] = dep_chan_vld_22_23;
    assign in_chan_dep_data_vec_23[25 : 0] = dep_chan_data_22_23;
    assign token_in_vec_23[0] = token_22_23;
    assign in_chan_dep_vld_vec_23[1] = dep_chan_vld_24_23;
    assign in_chan_dep_data_vec_23[51 : 26] = dep_chan_data_24_23;
    assign token_in_vec_23[1] = token_24_23;
    assign dep_chan_vld_23_22 = out_chan_dep_vld_vec_23[0];
    assign dep_chan_data_23_22 = out_chan_dep_data_23;
    assign token_23_22 = token_out_vec_23[0];
    assign dep_chan_vld_23_24 = out_chan_dep_vld_vec_23[1];
    assign dep_chan_data_23_24 = out_chan_dep_data_23;
    assign token_23_24 = token_out_vec_23[1];

    // Process: myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0
    alveo_hls4ml_hls_deadlock_detect_unit #(26, 24, 2, 2) alveo_hls4ml_hls_deadlock_detect_unit_24 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_24),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_24),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_24),
        .token_in_vec(token_in_vec_24),
        .dl_detect_in(dl_detect_out),
        .origin(origin[24]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_24),
        .out_chan_dep_data(out_chan_dep_data_24),
        .token_out_vec(token_out_vec_24),
        .dl_detect_out(dl_in_vec[24]));

    assign proc_24_data_FIFO_blk[0] = 1'b0 | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.layer23_out_0_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.layer23_out_1_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.layer23_out_2_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.layer23_out_3_blk_n);
    assign proc_24_data_PIPO_blk[0] = 1'b0;
    assign proc_24_start_FIFO_blk[0] = 1'b0 | (~myproject_U0.start_for_pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0_U.if_empty_n & myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.ap_idle & ~myproject_U0.start_for_pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0_U.if_write);
    assign proc_24_TLF_FIFO_blk[0] = 1'b0;
    assign proc_24_input_sync_blk[0] = 1'b0;
    assign proc_24_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_24[0] = dl_detect_out ? proc_dep_vld_vec_24_reg[0] : (proc_24_data_FIFO_blk[0] | proc_24_data_PIPO_blk[0] | proc_24_start_FIFO_blk[0] | proc_24_TLF_FIFO_blk[0] | proc_24_input_sync_blk[0] | proc_24_output_sync_blk[0]);
    assign proc_24_data_FIFO_blk[1] = 1'b0 | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_0_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_1_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_2_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_3_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_4_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_5_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_6_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_7_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_8_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_9_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_10_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_11_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_12_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_13_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_14_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_15_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_16_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_17_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_18_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_19_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_20_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_21_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_22_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_23_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_24_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_25_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_26_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_27_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_28_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_29_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_30_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_31_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_32_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_33_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_34_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_35_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_36_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_37_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_38_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_39_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_40_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_41_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_42_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_43_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_44_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_45_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_46_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_47_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_48_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_49_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_50_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_51_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_52_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_53_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_54_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_55_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_56_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_57_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_58_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_59_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_60_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_61_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_62_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_63_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_64_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_65_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_66_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_67_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_68_blk_n) | (~myproject_U0.pointwise_conv_1d_cl_ap_fixed_ap_fixed_16_6_5_3_0_config27_U0.out_stream_69_blk_n);
    assign proc_24_data_PIPO_blk[1] = 1'b0;
    assign proc_24_start_FIFO_blk[1] = 1'b0;
    assign proc_24_TLF_FIFO_blk[1] = 1'b0;
    assign proc_24_input_sync_blk[1] = 1'b0;
    assign proc_24_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_24[1] = dl_detect_out ? proc_dep_vld_vec_24_reg[1] : (proc_24_data_FIFO_blk[1] | proc_24_data_PIPO_blk[1] | proc_24_start_FIFO_blk[1] | proc_24_TLF_FIFO_blk[1] | proc_24_input_sync_blk[1] | proc_24_output_sync_blk[1]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_24_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_24_reg <= proc_dep_vld_vec_24;
        end
    end
    assign in_chan_dep_vld_vec_24[0] = dep_chan_vld_23_24;
    assign in_chan_dep_data_vec_24[25 : 0] = dep_chan_data_23_24;
    assign token_in_vec_24[0] = token_23_24;
    assign in_chan_dep_vld_vec_24[1] = dep_chan_vld_25_24;
    assign in_chan_dep_data_vec_24[51 : 26] = dep_chan_data_25_24;
    assign token_in_vec_24[1] = token_25_24;
    assign dep_chan_vld_24_23 = out_chan_dep_vld_vec_24[0];
    assign dep_chan_data_24_23 = out_chan_dep_data_24;
    assign token_24_23 = token_out_vec_24[0];
    assign dep_chan_vld_24_25 = out_chan_dep_vld_vec_24[1];
    assign dep_chan_data_24_25 = out_chan_dep_data_24;
    assign token_24_25 = token_out_vec_24[1];

    // Process: Loop_VITIS_LOOP_93_5_proc41_U0
    alveo_hls4ml_hls_deadlock_detect_unit #(26, 25, 3, 3) alveo_hls4ml_hls_deadlock_detect_unit_25 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_25),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_25),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_25),
        .token_in_vec(token_in_vec_25),
        .dl_detect_in(dl_detect_out),
        .origin(origin[25]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_25),
        .out_chan_dep_data(out_chan_dep_data_25),
        .token_out_vec(token_out_vec_25),
        .dl_detect_out(dl_in_vec[25]));

    assign proc_25_data_FIFO_blk[0] = 1'b0 | (~Loop_VITIS_LOOP_93_5_proc41_U0.out_r_blk_n);
    assign proc_25_data_PIPO_blk[0] = 1'b0;
    assign proc_25_start_FIFO_blk[0] = 1'b0 | (~start_for_Loop_VITIS_LOOP_93_5_proc41_U0_U.if_empty_n & Loop_VITIS_LOOP_93_5_proc41_U0.ap_idle & ~start_for_Loop_VITIS_LOOP_93_5_proc41_U0_U.if_write);
    assign proc_25_TLF_FIFO_blk[0] = 1'b0;
    assign proc_25_input_sync_blk[0] = 1'b0;
    assign proc_25_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_25[0] = dl_detect_out ? proc_dep_vld_vec_25_reg[0] : (proc_25_data_FIFO_blk[0] | proc_25_data_PIPO_blk[0] | proc_25_start_FIFO_blk[0] | proc_25_TLF_FIFO_blk[0] | proc_25_input_sync_blk[0] | proc_25_output_sync_blk[0]);
    assign proc_25_data_FIFO_blk[1] = 1'b0 | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_0_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_1_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_2_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_3_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_4_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_5_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_6_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_7_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_8_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_9_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_10_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_11_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_12_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_13_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_14_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_15_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_16_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_17_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_18_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_19_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_20_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_21_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_22_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_23_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_24_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_25_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_26_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_27_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_28_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_29_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_30_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_31_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_32_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_33_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_34_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_35_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_36_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_37_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_38_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_39_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_40_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_41_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_42_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_43_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_44_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_45_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_46_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_47_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_48_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_49_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_50_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_51_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_52_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_53_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_54_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_55_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_56_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_57_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_58_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_59_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_60_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_61_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_62_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_63_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_64_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_65_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_66_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_67_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_68_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_69_blk_n);
    assign proc_25_data_PIPO_blk[1] = 1'b0;
    assign proc_25_start_FIFO_blk[1] = 1'b0;
    assign proc_25_TLF_FIFO_blk[1] = 1'b0;
    assign proc_25_input_sync_blk[1] = 1'b0;
    assign proc_25_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_25[1] = dl_detect_out ? proc_dep_vld_vec_25_reg[1] : (proc_25_data_FIFO_blk[1] | proc_25_data_PIPO_blk[1] | proc_25_start_FIFO_blk[1] | proc_25_TLF_FIFO_blk[1] | proc_25_input_sync_blk[1] | proc_25_output_sync_blk[1]);
    assign proc_25_data_FIFO_blk[2] = 1'b0 | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_0_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_1_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_2_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_3_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_4_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_5_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_6_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_7_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_8_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_9_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_10_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_11_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_12_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_13_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_14_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_15_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_16_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_17_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_18_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_19_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_20_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_21_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_22_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_23_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_24_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_25_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_26_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_27_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_28_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_29_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_30_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_31_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_32_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_33_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_34_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_35_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_36_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_37_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_38_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_39_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_40_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_41_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_42_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_43_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_44_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_45_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_46_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_47_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_48_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_49_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_50_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_51_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_52_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_53_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_54_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_55_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_56_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_57_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_58_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_59_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_60_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_61_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_62_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_63_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_64_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_65_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_66_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_67_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_68_blk_n) | (~Loop_VITIS_LOOP_93_5_proc41_U0.grp_Loop_VITIS_LOOP_93_5_proc41_Pipeline_VITIS_LOOP_93_5_VITIS_LOOP_94_6_fu_202.out_stream_69_blk_n);
    assign proc_25_data_PIPO_blk[2] = 1'b0;
    assign proc_25_start_FIFO_blk[2] = 1'b0;
    assign proc_25_TLF_FIFO_blk[2] = 1'b0;
    assign proc_25_input_sync_blk[2] = 1'b0;
    assign proc_25_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_25[2] = dl_detect_out ? proc_dep_vld_vec_25_reg[2] : (proc_25_data_FIFO_blk[2] | proc_25_data_PIPO_blk[2] | proc_25_start_FIFO_blk[2] | proc_25_TLF_FIFO_blk[2] | proc_25_input_sync_blk[2] | proc_25_output_sync_blk[2]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_25_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_25_reg <= proc_dep_vld_vec_25;
        end
    end
    assign in_chan_dep_vld_vec_25[0] = dep_chan_vld_0_25;
    assign in_chan_dep_data_vec_25[25 : 0] = dep_chan_data_0_25;
    assign token_in_vec_25[0] = token_0_25;
    assign in_chan_dep_vld_vec_25[1] = dep_chan_vld_3_25;
    assign in_chan_dep_data_vec_25[51 : 26] = dep_chan_data_3_25;
    assign token_in_vec_25[1] = token_3_25;
    assign in_chan_dep_vld_vec_25[2] = dep_chan_vld_24_25;
    assign in_chan_dep_data_vec_25[77 : 52] = dep_chan_data_24_25;
    assign token_in_vec_25[2] = token_24_25;
    assign dep_chan_vld_25_0 = out_chan_dep_vld_vec_25[0];
    assign dep_chan_data_25_0 = out_chan_dep_data_25;
    assign token_25_0 = token_out_vec_25[0];
    assign dep_chan_vld_25_3 = out_chan_dep_vld_vec_25[1];
    assign dep_chan_data_25_3 = out_chan_dep_data_25;
    assign token_25_3 = token_out_vec_25[1];
    assign dep_chan_vld_25_24 = out_chan_dep_vld_vec_25[2];
    assign dep_chan_data_25_24 = out_chan_dep_data_25;
    assign token_25_24 = token_out_vec_25[2];


`include "alveo_hls4ml_hls_deadlock_report_unit.vh"
